`timescale 1 ns / 1 ps

module AESL_deadlock_detector (
    input dl_reset,
    input all_finish,
    input dl_clock);

    wire [6:0] proc_0_data_FIFO_blk;
    wire [6:0] proc_0_data_PIPO_blk;
    wire [6:0] proc_0_start_FIFO_blk;
    wire [6:0] proc_0_TLF_FIFO_blk;
    wire [6:0] proc_0_input_sync_blk;
    wire [6:0] proc_0_output_sync_blk;
    wire [6:0] proc_dep_vld_vec_0;
    reg [6:0] proc_dep_vld_vec_0_reg;
    wire [6:0] in_chan_dep_vld_vec_0;
    wire [118:0] in_chan_dep_data_vec_0;
    wire [6:0] token_in_vec_0;
    wire [6:0] out_chan_dep_vld_vec_0;
    wire [16:0] out_chan_dep_data_0;
    wire [6:0] token_out_vec_0;
    wire dl_detect_out_0;
    wire dep_chan_vld_1_0;
    wire [16:0] dep_chan_data_1_0;
    wire token_1_0;
    wire dep_chan_vld_2_0;
    wire [16:0] dep_chan_data_2_0;
    wire token_2_0;
    wire dep_chan_vld_3_0;
    wire [16:0] dep_chan_data_3_0;
    wire token_3_0;
    wire dep_chan_vld_4_0;
    wire [16:0] dep_chan_data_4_0;
    wire token_4_0;
    wire dep_chan_vld_5_0;
    wire [16:0] dep_chan_data_5_0;
    wire token_5_0;
    wire dep_chan_vld_7_0;
    wire [16:0] dep_chan_data_7_0;
    wire token_7_0;
    wire dep_chan_vld_16_0;
    wire [16:0] dep_chan_data_16_0;
    wire token_16_0;
    wire [3:0] proc_1_data_FIFO_blk;
    wire [3:0] proc_1_data_PIPO_blk;
    wire [3:0] proc_1_start_FIFO_blk;
    wire [3:0] proc_1_TLF_FIFO_blk;
    wire [3:0] proc_1_input_sync_blk;
    wire [3:0] proc_1_output_sync_blk;
    wire [3:0] proc_dep_vld_vec_1;
    reg [3:0] proc_dep_vld_vec_1_reg;
    wire [8:0] in_chan_dep_vld_vec_1;
    wire [152:0] in_chan_dep_data_vec_1;
    wire [8:0] token_in_vec_1;
    wire [3:0] out_chan_dep_vld_vec_1;
    wire [16:0] out_chan_dep_data_1;
    wire [3:0] token_out_vec_1;
    wire dl_detect_out_1;
    wire dep_chan_vld_0_1;
    wire [16:0] dep_chan_data_0_1;
    wire token_0_1;
    wire dep_chan_vld_2_1;
    wire [16:0] dep_chan_data_2_1;
    wire token_2_1;
    wire dep_chan_vld_3_1;
    wire [16:0] dep_chan_data_3_1;
    wire token_3_1;
    wire dep_chan_vld_6_1;
    wire [16:0] dep_chan_data_6_1;
    wire token_6_1;
    wire dep_chan_vld_7_1;
    wire [16:0] dep_chan_data_7_1;
    wire token_7_1;
    wire dep_chan_vld_8_1;
    wire [16:0] dep_chan_data_8_1;
    wire token_8_1;
    wire dep_chan_vld_9_1;
    wire [16:0] dep_chan_data_9_1;
    wire token_9_1;
    wire dep_chan_vld_11_1;
    wire [16:0] dep_chan_data_11_1;
    wire token_11_1;
    wire dep_chan_vld_13_1;
    wire [16:0] dep_chan_data_13_1;
    wire token_13_1;
    wire [5:0] proc_2_data_FIFO_blk;
    wire [5:0] proc_2_data_PIPO_blk;
    wire [5:0] proc_2_start_FIFO_blk;
    wire [5:0] proc_2_TLF_FIFO_blk;
    wire [5:0] proc_2_input_sync_blk;
    wire [5:0] proc_2_output_sync_blk;
    wire [5:0] proc_dep_vld_vec_2;
    reg [5:0] proc_dep_vld_vec_2_reg;
    wire [5:0] in_chan_dep_vld_vec_2;
    wire [101:0] in_chan_dep_data_vec_2;
    wire [5:0] token_in_vec_2;
    wire [5:0] out_chan_dep_vld_vec_2;
    wire [16:0] out_chan_dep_data_2;
    wire [5:0] token_out_vec_2;
    wire dl_detect_out_2;
    wire dep_chan_vld_0_2;
    wire [16:0] dep_chan_data_0_2;
    wire token_0_2;
    wire dep_chan_vld_1_2;
    wire [16:0] dep_chan_data_1_2;
    wire token_1_2;
    wire dep_chan_vld_3_2;
    wire [16:0] dep_chan_data_3_2;
    wire token_3_2;
    wire dep_chan_vld_7_2;
    wire [16:0] dep_chan_data_7_2;
    wire token_7_2;
    wire dep_chan_vld_14_2;
    wire [16:0] dep_chan_data_14_2;
    wire token_14_2;
    wire dep_chan_vld_15_2;
    wire [16:0] dep_chan_data_15_2;
    wire token_15_2;
    wire [5:0] proc_3_data_FIFO_blk;
    wire [5:0] proc_3_data_PIPO_blk;
    wire [5:0] proc_3_start_FIFO_blk;
    wire [5:0] proc_3_TLF_FIFO_blk;
    wire [5:0] proc_3_input_sync_blk;
    wire [5:0] proc_3_output_sync_blk;
    wire [5:0] proc_dep_vld_vec_3;
    reg [5:0] proc_dep_vld_vec_3_reg;
    wire [5:0] in_chan_dep_vld_vec_3;
    wire [101:0] in_chan_dep_data_vec_3;
    wire [5:0] token_in_vec_3;
    wire [5:0] out_chan_dep_vld_vec_3;
    wire [16:0] out_chan_dep_data_3;
    wire [5:0] token_out_vec_3;
    wire dl_detect_out_3;
    wire dep_chan_vld_0_3;
    wire [16:0] dep_chan_data_0_3;
    wire token_0_3;
    wire dep_chan_vld_1_3;
    wire [16:0] dep_chan_data_1_3;
    wire token_1_3;
    wire dep_chan_vld_2_3;
    wire [16:0] dep_chan_data_2_3;
    wire token_2_3;
    wire dep_chan_vld_4_3;
    wire [16:0] dep_chan_data_4_3;
    wire token_4_3;
    wire dep_chan_vld_6_3;
    wire [16:0] dep_chan_data_6_3;
    wire token_6_3;
    wire dep_chan_vld_7_3;
    wire [16:0] dep_chan_data_7_3;
    wire token_7_3;
    wire [2:0] proc_4_data_FIFO_blk;
    wire [2:0] proc_4_data_PIPO_blk;
    wire [2:0] proc_4_start_FIFO_blk;
    wire [2:0] proc_4_TLF_FIFO_blk;
    wire [2:0] proc_4_input_sync_blk;
    wire [2:0] proc_4_output_sync_blk;
    wire [2:0] proc_dep_vld_vec_4;
    reg [2:0] proc_dep_vld_vec_4_reg;
    wire [2:0] in_chan_dep_vld_vec_4;
    wire [50:0] in_chan_dep_data_vec_4;
    wire [2:0] token_in_vec_4;
    wire [2:0] out_chan_dep_vld_vec_4;
    wire [16:0] out_chan_dep_data_4;
    wire [2:0] token_out_vec_4;
    wire dl_detect_out_4;
    wire dep_chan_vld_0_4;
    wire [16:0] dep_chan_data_0_4;
    wire token_0_4;
    wire dep_chan_vld_3_4;
    wire [16:0] dep_chan_data_3_4;
    wire token_3_4;
    wire dep_chan_vld_5_4;
    wire [16:0] dep_chan_data_5_4;
    wire token_5_4;
    wire [5:0] proc_5_data_FIFO_blk;
    wire [5:0] proc_5_data_PIPO_blk;
    wire [5:0] proc_5_start_FIFO_blk;
    wire [5:0] proc_5_TLF_FIFO_blk;
    wire [5:0] proc_5_input_sync_blk;
    wire [5:0] proc_5_output_sync_blk;
    wire [5:0] proc_dep_vld_vec_5;
    reg [5:0] proc_dep_vld_vec_5_reg;
    wire [5:0] in_chan_dep_vld_vec_5;
    wire [101:0] in_chan_dep_data_vec_5;
    wire [5:0] token_in_vec_5;
    wire [5:0] out_chan_dep_vld_vec_5;
    wire [16:0] out_chan_dep_data_5;
    wire [5:0] token_out_vec_5;
    wire dl_detect_out_5;
    wire dep_chan_vld_0_5;
    wire [16:0] dep_chan_data_0_5;
    wire token_0_5;
    wire dep_chan_vld_4_5;
    wire [16:0] dep_chan_data_4_5;
    wire token_4_5;
    wire dep_chan_vld_6_5;
    wire [16:0] dep_chan_data_6_5;
    wire token_6_5;
    wire dep_chan_vld_12_5;
    wire [16:0] dep_chan_data_12_5;
    wire token_12_5;
    wire dep_chan_vld_13_5;
    wire [16:0] dep_chan_data_13_5;
    wire token_13_5;
    wire dep_chan_vld_16_5;
    wire [16:0] dep_chan_data_16_5;
    wire token_16_5;
    wire [3:0] proc_6_data_FIFO_blk;
    wire [3:0] proc_6_data_PIPO_blk;
    wire [3:0] proc_6_start_FIFO_blk;
    wire [3:0] proc_6_TLF_FIFO_blk;
    wire [3:0] proc_6_input_sync_blk;
    wire [3:0] proc_6_output_sync_blk;
    wire [3:0] proc_dep_vld_vec_6;
    reg [3:0] proc_dep_vld_vec_6_reg;
    wire [2:0] in_chan_dep_vld_vec_6;
    wire [50:0] in_chan_dep_data_vec_6;
    wire [2:0] token_in_vec_6;
    wire [3:0] out_chan_dep_vld_vec_6;
    wire [16:0] out_chan_dep_data_6;
    wire [3:0] token_out_vec_6;
    wire dl_detect_out_6;
    wire dep_chan_vld_3_6;
    wire [16:0] dep_chan_data_3_6;
    wire token_3_6;
    wire dep_chan_vld_5_6;
    wire [16:0] dep_chan_data_5_6;
    wire token_5_6;
    wire dep_chan_vld_11_6;
    wire [16:0] dep_chan_data_11_6;
    wire token_11_6;
    wire [5:0] proc_7_data_FIFO_blk;
    wire [5:0] proc_7_data_PIPO_blk;
    wire [5:0] proc_7_start_FIFO_blk;
    wire [5:0] proc_7_TLF_FIFO_blk;
    wire [5:0] proc_7_input_sync_blk;
    wire [5:0] proc_7_output_sync_blk;
    wire [5:0] proc_dep_vld_vec_7;
    reg [5:0] proc_dep_vld_vec_7_reg;
    wire [5:0] in_chan_dep_vld_vec_7;
    wire [101:0] in_chan_dep_data_vec_7;
    wire [5:0] token_in_vec_7;
    wire [5:0] out_chan_dep_vld_vec_7;
    wire [16:0] out_chan_dep_data_7;
    wire [5:0] token_out_vec_7;
    wire dl_detect_out_7;
    wire dep_chan_vld_0_7;
    wire [16:0] dep_chan_data_0_7;
    wire token_0_7;
    wire dep_chan_vld_1_7;
    wire [16:0] dep_chan_data_1_7;
    wire token_1_7;
    wire dep_chan_vld_2_7;
    wire [16:0] dep_chan_data_2_7;
    wire token_2_7;
    wire dep_chan_vld_3_7;
    wire [16:0] dep_chan_data_3_7;
    wire token_3_7;
    wire dep_chan_vld_8_7;
    wire [16:0] dep_chan_data_8_7;
    wire token_8_7;
    wire dep_chan_vld_9_7;
    wire [16:0] dep_chan_data_9_7;
    wire token_9_7;
    wire [2:0] proc_8_data_FIFO_blk;
    wire [2:0] proc_8_data_PIPO_blk;
    wire [2:0] proc_8_start_FIFO_blk;
    wire [2:0] proc_8_TLF_FIFO_blk;
    wire [2:0] proc_8_input_sync_blk;
    wire [2:0] proc_8_output_sync_blk;
    wire [2:0] proc_dep_vld_vec_8;
    reg [2:0] proc_dep_vld_vec_8_reg;
    wire [1:0] in_chan_dep_vld_vec_8;
    wire [33:0] in_chan_dep_data_vec_8;
    wire [1:0] token_in_vec_8;
    wire [2:0] out_chan_dep_vld_vec_8;
    wire [16:0] out_chan_dep_data_8;
    wire [2:0] token_out_vec_8;
    wire dl_detect_out_8;
    wire dep_chan_vld_7_8;
    wire [16:0] dep_chan_data_7_8;
    wire token_7_8;
    wire dep_chan_vld_10_8;
    wire [16:0] dep_chan_data_10_8;
    wire token_10_8;
    wire [2:0] proc_9_data_FIFO_blk;
    wire [2:0] proc_9_data_PIPO_blk;
    wire [2:0] proc_9_start_FIFO_blk;
    wire [2:0] proc_9_TLF_FIFO_blk;
    wire [2:0] proc_9_input_sync_blk;
    wire [2:0] proc_9_output_sync_blk;
    wire [2:0] proc_dep_vld_vec_9;
    reg [2:0] proc_dep_vld_vec_9_reg;
    wire [1:0] in_chan_dep_vld_vec_9;
    wire [33:0] in_chan_dep_data_vec_9;
    wire [1:0] token_in_vec_9;
    wire [2:0] out_chan_dep_vld_vec_9;
    wire [16:0] out_chan_dep_data_9;
    wire [2:0] token_out_vec_9;
    wire dl_detect_out_9;
    wire dep_chan_vld_7_9;
    wire [16:0] dep_chan_data_7_9;
    wire token_7_9;
    wire dep_chan_vld_10_9;
    wire [16:0] dep_chan_data_10_9;
    wire token_10_9;
    wire [2:0] proc_10_data_FIFO_blk;
    wire [2:0] proc_10_data_PIPO_blk;
    wire [2:0] proc_10_start_FIFO_blk;
    wire [2:0] proc_10_TLF_FIFO_blk;
    wire [2:0] proc_10_input_sync_blk;
    wire [2:0] proc_10_output_sync_blk;
    wire [2:0] proc_dep_vld_vec_10;
    reg [2:0] proc_dep_vld_vec_10_reg;
    wire [2:0] in_chan_dep_vld_vec_10;
    wire [50:0] in_chan_dep_data_vec_10;
    wire [2:0] token_in_vec_10;
    wire [2:0] out_chan_dep_vld_vec_10;
    wire [16:0] out_chan_dep_data_10;
    wire [2:0] token_out_vec_10;
    wire dl_detect_out_10;
    wire dep_chan_vld_8_10;
    wire [16:0] dep_chan_data_8_10;
    wire token_8_10;
    wire dep_chan_vld_9_10;
    wire [16:0] dep_chan_data_9_10;
    wire token_9_10;
    wire dep_chan_vld_11_10;
    wire [16:0] dep_chan_data_11_10;
    wire token_11_10;
    wire [4:0] proc_11_data_FIFO_blk;
    wire [4:0] proc_11_data_PIPO_blk;
    wire [4:0] proc_11_start_FIFO_blk;
    wire [4:0] proc_11_TLF_FIFO_blk;
    wire [4:0] proc_11_input_sync_blk;
    wire [4:0] proc_11_output_sync_blk;
    wire [4:0] proc_dep_vld_vec_11;
    reg [4:0] proc_dep_vld_vec_11_reg;
    wire [3:0] in_chan_dep_vld_vec_11;
    wire [67:0] in_chan_dep_data_vec_11;
    wire [3:0] token_in_vec_11;
    wire [4:0] out_chan_dep_vld_vec_11;
    wire [16:0] out_chan_dep_data_11;
    wire [4:0] token_out_vec_11;
    wire dl_detect_out_11;
    wire dep_chan_vld_6_11;
    wire [16:0] dep_chan_data_6_11;
    wire token_6_11;
    wire dep_chan_vld_10_11;
    wire [16:0] dep_chan_data_10_11;
    wire token_10_11;
    wire dep_chan_vld_12_11;
    wire [16:0] dep_chan_data_12_11;
    wire token_12_11;
    wire dep_chan_vld_13_11;
    wire [16:0] dep_chan_data_13_11;
    wire token_13_11;
    wire [3:0] proc_12_data_FIFO_blk;
    wire [3:0] proc_12_data_PIPO_blk;
    wire [3:0] proc_12_start_FIFO_blk;
    wire [3:0] proc_12_TLF_FIFO_blk;
    wire [3:0] proc_12_input_sync_blk;
    wire [3:0] proc_12_output_sync_blk;
    wire [3:0] proc_dep_vld_vec_12;
    reg [3:0] proc_dep_vld_vec_12_reg;
    wire [3:0] in_chan_dep_vld_vec_12;
    wire [67:0] in_chan_dep_data_vec_12;
    wire [3:0] token_in_vec_12;
    wire [3:0] out_chan_dep_vld_vec_12;
    wire [16:0] out_chan_dep_data_12;
    wire [3:0] token_out_vec_12;
    wire dl_detect_out_12;
    wire dep_chan_vld_5_12;
    wire [16:0] dep_chan_data_5_12;
    wire token_5_12;
    wire dep_chan_vld_11_12;
    wire [16:0] dep_chan_data_11_12;
    wire token_11_12;
    wire dep_chan_vld_13_12;
    wire [16:0] dep_chan_data_13_12;
    wire token_13_12;
    wire dep_chan_vld_16_12;
    wire [16:0] dep_chan_data_16_12;
    wire token_16_12;
    wire [5:0] proc_13_data_FIFO_blk;
    wire [5:0] proc_13_data_PIPO_blk;
    wire [5:0] proc_13_start_FIFO_blk;
    wire [5:0] proc_13_TLF_FIFO_blk;
    wire [5:0] proc_13_input_sync_blk;
    wire [5:0] proc_13_output_sync_blk;
    wire [5:0] proc_dep_vld_vec_13;
    reg [5:0] proc_dep_vld_vec_13_reg;
    wire [4:0] in_chan_dep_vld_vec_13;
    wire [84:0] in_chan_dep_data_vec_13;
    wire [4:0] token_in_vec_13;
    wire [5:0] out_chan_dep_vld_vec_13;
    wire [16:0] out_chan_dep_data_13;
    wire [5:0] token_out_vec_13;
    wire dl_detect_out_13;
    wire dep_chan_vld_5_13;
    wire [16:0] dep_chan_data_5_13;
    wire token_5_13;
    wire dep_chan_vld_11_13;
    wire [16:0] dep_chan_data_11_13;
    wire token_11_13;
    wire dep_chan_vld_12_13;
    wire [16:0] dep_chan_data_12_13;
    wire token_12_13;
    wire dep_chan_vld_14_13;
    wire [16:0] dep_chan_data_14_13;
    wire token_14_13;
    wire dep_chan_vld_16_13;
    wire [16:0] dep_chan_data_16_13;
    wire token_16_13;
    wire [2:0] proc_14_data_FIFO_blk;
    wire [2:0] proc_14_data_PIPO_blk;
    wire [2:0] proc_14_start_FIFO_blk;
    wire [2:0] proc_14_TLF_FIFO_blk;
    wire [2:0] proc_14_input_sync_blk;
    wire [2:0] proc_14_output_sync_blk;
    wire [2:0] proc_dep_vld_vec_14;
    reg [2:0] proc_dep_vld_vec_14_reg;
    wire [2:0] in_chan_dep_vld_vec_14;
    wire [50:0] in_chan_dep_data_vec_14;
    wire [2:0] token_in_vec_14;
    wire [2:0] out_chan_dep_vld_vec_14;
    wire [16:0] out_chan_dep_data_14;
    wire [2:0] token_out_vec_14;
    wire dl_detect_out_14;
    wire dep_chan_vld_2_14;
    wire [16:0] dep_chan_data_2_14;
    wire token_2_14;
    wire dep_chan_vld_13_14;
    wire [16:0] dep_chan_data_13_14;
    wire token_13_14;
    wire dep_chan_vld_15_14;
    wire [16:0] dep_chan_data_15_14;
    wire token_15_14;
    wire [2:0] proc_15_data_FIFO_blk;
    wire [2:0] proc_15_data_PIPO_blk;
    wire [2:0] proc_15_start_FIFO_blk;
    wire [2:0] proc_15_TLF_FIFO_blk;
    wire [2:0] proc_15_input_sync_blk;
    wire [2:0] proc_15_output_sync_blk;
    wire [2:0] proc_dep_vld_vec_15;
    reg [2:0] proc_dep_vld_vec_15_reg;
    wire [2:0] in_chan_dep_vld_vec_15;
    wire [50:0] in_chan_dep_data_vec_15;
    wire [2:0] token_in_vec_15;
    wire [2:0] out_chan_dep_vld_vec_15;
    wire [16:0] out_chan_dep_data_15;
    wire [2:0] token_out_vec_15;
    wire dl_detect_out_15;
    wire dep_chan_vld_2_15;
    wire [16:0] dep_chan_data_2_15;
    wire token_2_15;
    wire dep_chan_vld_14_15;
    wire [16:0] dep_chan_data_14_15;
    wire token_14_15;
    wire dep_chan_vld_16_15;
    wire [16:0] dep_chan_data_16_15;
    wire token_16_15;
    wire [4:0] proc_16_data_FIFO_blk;
    wire [4:0] proc_16_data_PIPO_blk;
    wire [4:0] proc_16_start_FIFO_blk;
    wire [4:0] proc_16_TLF_FIFO_blk;
    wire [4:0] proc_16_input_sync_blk;
    wire [4:0] proc_16_output_sync_blk;
    wire [4:0] proc_dep_vld_vec_16;
    reg [4:0] proc_dep_vld_vec_16_reg;
    wire [4:0] in_chan_dep_vld_vec_16;
    wire [84:0] in_chan_dep_data_vec_16;
    wire [4:0] token_in_vec_16;
    wire [4:0] out_chan_dep_vld_vec_16;
    wire [16:0] out_chan_dep_data_16;
    wire [4:0] token_out_vec_16;
    wire dl_detect_out_16;
    wire dep_chan_vld_0_16;
    wire [16:0] dep_chan_data_0_16;
    wire token_0_16;
    wire dep_chan_vld_5_16;
    wire [16:0] dep_chan_data_5_16;
    wire token_5_16;
    wire dep_chan_vld_12_16;
    wire [16:0] dep_chan_data_12_16;
    wire token_12_16;
    wire dep_chan_vld_13_16;
    wire [16:0] dep_chan_data_13_16;
    wire token_13_16;
    wire dep_chan_vld_15_16;
    wire [16:0] dep_chan_data_15_16;
    wire token_15_16;
    wire [16:0] dl_in_vec;
    wire dl_detect_out;
    wire token_clear;
    wire [16:0] origin;

    reg ap_done_reg_0;// for module AESL_inst_top.ConvertInputToArray_U0
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            ap_done_reg_0 <= 'b0;
        end
        else begin
            ap_done_reg_0 <= AESL_inst_top.ConvertInputToArray_U0.ap_done & ~AESL_inst_top.ConvertInputToArray_U0.ap_continue;
        end
    end

    reg ap_done_reg_1;// for module AESL_inst_top.ConvWeightToArray_U0
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            ap_done_reg_1 <= 'b0;
        end
        else begin
            ap_done_reg_1 <= AESL_inst_top.ConvWeightToArray_U0.ap_done & ~AESL_inst_top.ConvWeightToArray_U0.ap_continue;
        end
    end

    reg ap_done_reg_2;// for module AESL_inst_top.MMWeightToArray_U0
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            ap_done_reg_2 <= 'b0;
        end
        else begin
            ap_done_reg_2 <= AESL_inst_top.MMWeightToArray_U0.ap_done & ~AESL_inst_top.MMWeightToArray_U0.ap_continue;
        end
    end

    reg ap_done_reg_3;// for module AESL_inst_top.Compute_U0
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            ap_done_reg_3 <= 'b0;
        end
        else begin
            ap_done_reg_3 <= AESL_inst_top.Compute_U0.ap_done & ~AESL_inst_top.Compute_U0.ap_continue;
        end
    end

    reg ap_done_reg_4;// for module AESL_inst_top.ConvToOutStream_U0
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            ap_done_reg_4 <= 'b0;
        end
        else begin
            ap_done_reg_4 <= AESL_inst_top.ConvToOutStream_U0.ap_done & ~AESL_inst_top.ConvToOutStream_U0.ap_continue;
        end
    end

reg [15:0] trans_in_cnt_0;// for process AESL_inst_top.entry_proc_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_0 <= 16'h0;
    end
    else if (AESL_inst_top.entry_proc_U0.start_write == 1'b1) begin
        trans_in_cnt_0 <= trans_in_cnt_0 + 16'h1;
    end
    else begin
        trans_in_cnt_0 <= trans_in_cnt_0;
    end
end

reg [15:0] trans_out_cnt_0;// for process AESL_inst_top.entry_proc_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_0 <= 16'h0;
    end
    else if (AESL_inst_top.entry_proc_U0.ap_done == 1'b1 && AESL_inst_top.entry_proc_U0.ap_continue == 1'b1) begin
        trans_out_cnt_0 <= trans_out_cnt_0 + 16'h1;
    end
    else begin
        trans_out_cnt_0 <= trans_out_cnt_0;
    end
end

reg [15:0] trans_in_cnt_1;// for process AESL_inst_top.ConvWeightToArray_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_1 <= 16'h0;
    end
    else if (AESL_inst_top.ConvWeightToArray_U0.start_write == 1'b1) begin
        trans_in_cnt_1 <= trans_in_cnt_1 + 16'h1;
    end
    else begin
        trans_in_cnt_1 <= trans_in_cnt_1;
    end
end

reg [15:0] trans_out_cnt_1;// for process AESL_inst_top.ConvWeightToArray_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_1 <= 16'h0;
    end
    else if (AESL_inst_top.ConvWeightToArray_U0.ap_done == 1'b1 && AESL_inst_top.ConvWeightToArray_U0.ap_continue == 1'b1) begin
        trans_out_cnt_1 <= trans_out_cnt_1 + 16'h1;
    end
    else begin
        trans_out_cnt_1 <= trans_out_cnt_1;
    end
end

reg [15:0] trans_in_cnt_2;// for process AESL_inst_top.Sliding_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_2 <= 16'h0;
    end
    else if (AESL_inst_top.Sliding_U0.start_write == 1'b1) begin
        trans_in_cnt_2 <= trans_in_cnt_2 + 16'h1;
    end
    else begin
        trans_in_cnt_2 <= trans_in_cnt_2;
    end
end

reg [15:0] trans_out_cnt_2;// for process AESL_inst_top.Sliding_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_2 <= 16'h0;
    end
    else if (AESL_inst_top.Sliding_U0.ap_done == 1'b1 && AESL_inst_top.Sliding_U0.ap_continue == 1'b1) begin
        trans_out_cnt_2 <= trans_out_cnt_2 + 16'h1;
    end
    else begin
        trans_out_cnt_2 <= trans_out_cnt_2;
    end
end

reg [15:0] trans_in_cnt_3;// for process AESL_inst_top.ConvertBias_BN_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_3 <= 16'h0;
    end
    else if (AESL_inst_top.ConvertBias_BN_U0.start_write == 1'b1) begin
        trans_in_cnt_3 <= trans_in_cnt_3 + 16'h1;
    end
    else begin
        trans_in_cnt_3 <= trans_in_cnt_3;
    end
end

reg [15:0] trans_out_cnt_3;// for process AESL_inst_top.ConvertBias_BN_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_3 <= 16'h0;
    end
    else if (AESL_inst_top.ConvertBias_BN_U0.ap_done == 1'b1 && AESL_inst_top.ConvertBias_BN_U0.ap_continue == 1'b1) begin
        trans_out_cnt_3 <= trans_out_cnt_3 + 16'h1;
    end
    else begin
        trans_out_cnt_3 <= trans_out_cnt_3;
    end
end

    // Process: AESL_inst_top.entry_proc_U0
    AESL_deadlock_detect_unit #(17, 0, 7, 7) AESL_deadlock_detect_unit_0 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_0),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_0),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_0),
        .token_in_vec(token_in_vec_0),
        .dl_detect_in(dl_detect_out),
        .origin(origin[0]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_0),
        .out_chan_dep_data(out_chan_dep_data_0),
        .token_out_vec(token_out_vec_0),
        .dl_detect_out(dl_in_vec[0]));

    assign proc_0_data_FIFO_blk[0] = 1'b0 | (~AESL_inst_top.entry_proc_U0.Output_r_c_blk_n);
    assign proc_0_data_PIPO_blk[0] = 1'b0;
    assign proc_0_start_FIFO_blk[0] = 1'b0 | (~AESL_inst_top.start_for_ResOutput_U0_U.if_full_n & AESL_inst_top.entry_proc_U0.ap_start & ~AESL_inst_top.entry_proc_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~AESL_inst_top.start_for_ResOutput_U0_U.if_read);
    assign proc_0_TLF_FIFO_blk[0] = 1'b0;
    assign proc_0_input_sync_blk[0] = 1'b0;
    assign proc_0_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_0[0] = dl_detect_out ? proc_dep_vld_vec_0_reg[0] : (proc_0_data_FIFO_blk[0] | proc_0_data_PIPO_blk[0] | proc_0_start_FIFO_blk[0] | proc_0_TLF_FIFO_blk[0] | proc_0_input_sync_blk[0] | proc_0_output_sync_blk[0]);
    assign proc_0_data_FIFO_blk[1] = 1'b0 | (~AESL_inst_top.entry_proc_U0.K_c58_blk_n) | (~AESL_inst_top.entry_proc_U0.S_c61_blk_n);
    assign proc_0_data_PIPO_blk[1] = 1'b0;
    assign proc_0_start_FIFO_blk[1] = 1'b0 | (~AESL_inst_top.start_for_Sliding_U0_U.if_full_n & AESL_inst_top.entry_proc_U0.ap_start & ~AESL_inst_top.entry_proc_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~AESL_inst_top.start_for_Sliding_U0_U.if_read);
    assign proc_0_TLF_FIFO_blk[1] = 1'b0;
    assign proc_0_input_sync_blk[1] = 1'b0;
    assign proc_0_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_0[1] = dl_detect_out ? proc_dep_vld_vec_0_reg[1] : (proc_0_data_FIFO_blk[1] | proc_0_data_PIPO_blk[1] | proc_0_start_FIFO_blk[1] | proc_0_TLF_FIFO_blk[1] | proc_0_input_sync_blk[1] | proc_0_output_sync_blk[1]);
    assign proc_0_data_FIFO_blk[2] = 1'b0 | (~AESL_inst_top.entry_proc_U0.P_c60_blk_n);
    assign proc_0_data_PIPO_blk[2] = 1'b0;
    assign proc_0_start_FIFO_blk[2] = 1'b0 | (~AESL_inst_top.start_for_Padding_U0_U.if_full_n & AESL_inst_top.entry_proc_U0.ap_start & ~AESL_inst_top.entry_proc_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~AESL_inst_top.start_for_Padding_U0_U.if_read);
    assign proc_0_TLF_FIFO_blk[2] = 1'b0;
    assign proc_0_input_sync_blk[2] = 1'b0;
    assign proc_0_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_0[2] = dl_detect_out ? proc_dep_vld_vec_0_reg[2] : (proc_0_data_FIFO_blk[2] | proc_0_data_PIPO_blk[2] | proc_0_start_FIFO_blk[2] | proc_0_TLF_FIFO_blk[2] | proc_0_input_sync_blk[2] | proc_0_output_sync_blk[2]);
    assign proc_0_data_FIFO_blk[3] = 1'b0;
    assign proc_0_data_PIPO_blk[3] = 1'b0;
    assign proc_0_start_FIFO_blk[3] = 1'b0;
    assign proc_0_TLF_FIFO_blk[3] = 1'b0;
    assign proc_0_input_sync_blk[3] = 1'b0 | (AESL_inst_top.ap_sync_entry_proc_U0_ap_ready & AESL_inst_top.entry_proc_U0.ap_idle & ~AESL_inst_top.ap_sync_Block_entry3_proc_U0_ap_ready);
    assign proc_0_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_0[3] = dl_detect_out ? proc_dep_vld_vec_0_reg[3] : (proc_0_data_FIFO_blk[3] | proc_0_data_PIPO_blk[3] | proc_0_start_FIFO_blk[3] | proc_0_TLF_FIFO_blk[3] | proc_0_input_sync_blk[3] | proc_0_output_sync_blk[3]);
    assign proc_0_data_FIFO_blk[4] = 1'b0;
    assign proc_0_data_PIPO_blk[4] = 1'b0;
    assign proc_0_start_FIFO_blk[4] = 1'b0;
    assign proc_0_TLF_FIFO_blk[4] = 1'b0;
    assign proc_0_input_sync_blk[4] = 1'b0 | (AESL_inst_top.ap_sync_entry_proc_U0_ap_ready & AESL_inst_top.entry_proc_U0.ap_idle & ~AESL_inst_top.ap_sync_ConvertBias_BN_U0_ap_ready);
    assign proc_0_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_0[4] = dl_detect_out ? proc_dep_vld_vec_0_reg[4] : (proc_0_data_FIFO_blk[4] | proc_0_data_PIPO_blk[4] | proc_0_start_FIFO_blk[4] | proc_0_TLF_FIFO_blk[4] | proc_0_input_sync_blk[4] | proc_0_output_sync_blk[4]);
    assign proc_0_data_FIFO_blk[5] = 1'b0;
    assign proc_0_data_PIPO_blk[5] = 1'b0;
    assign proc_0_start_FIFO_blk[5] = 1'b0;
    assign proc_0_TLF_FIFO_blk[5] = 1'b0;
    assign proc_0_input_sync_blk[5] = 1'b0 | (AESL_inst_top.ap_sync_entry_proc_U0_ap_ready & AESL_inst_top.entry_proc_U0.ap_idle & ~AESL_inst_top.ap_sync_ConvertInputToStream_U0_ap_ready);
    assign proc_0_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_0[5] = dl_detect_out ? proc_dep_vld_vec_0_reg[5] : (proc_0_data_FIFO_blk[5] | proc_0_data_PIPO_blk[5] | proc_0_start_FIFO_blk[5] | proc_0_TLF_FIFO_blk[5] | proc_0_input_sync_blk[5] | proc_0_output_sync_blk[5]);
    assign proc_0_data_FIFO_blk[6] = 1'b0;
    assign proc_0_data_PIPO_blk[6] = 1'b0;
    assign proc_0_start_FIFO_blk[6] = 1'b0;
    assign proc_0_TLF_FIFO_blk[6] = 1'b0;
    assign proc_0_input_sync_blk[6] = 1'b0 | (AESL_inst_top.ap_sync_entry_proc_U0_ap_ready & AESL_inst_top.entry_proc_U0.ap_idle & ~AESL_inst_top.ap_sync_ConvertWeightToStream_U0_ap_ready);
    assign proc_0_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_0[6] = dl_detect_out ? proc_dep_vld_vec_0_reg[6] : (proc_0_data_FIFO_blk[6] | proc_0_data_PIPO_blk[6] | proc_0_start_FIFO_blk[6] | proc_0_TLF_FIFO_blk[6] | proc_0_input_sync_blk[6] | proc_0_output_sync_blk[6]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_0_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_0_reg <= proc_dep_vld_vec_0;
        end
    end
    assign in_chan_dep_vld_vec_0[0] = dep_chan_vld_1_0;
    assign in_chan_dep_data_vec_0[16 : 0] = dep_chan_data_1_0;
    assign token_in_vec_0[0] = token_1_0;
    assign in_chan_dep_vld_vec_0[1] = dep_chan_vld_2_0;
    assign in_chan_dep_data_vec_0[33 : 17] = dep_chan_data_2_0;
    assign token_in_vec_0[1] = token_2_0;
    assign in_chan_dep_vld_vec_0[2] = dep_chan_vld_3_0;
    assign in_chan_dep_data_vec_0[50 : 34] = dep_chan_data_3_0;
    assign token_in_vec_0[2] = token_3_0;
    assign in_chan_dep_vld_vec_0[3] = dep_chan_vld_4_0;
    assign in_chan_dep_data_vec_0[67 : 51] = dep_chan_data_4_0;
    assign token_in_vec_0[3] = token_4_0;
    assign in_chan_dep_vld_vec_0[4] = dep_chan_vld_5_0;
    assign in_chan_dep_data_vec_0[84 : 68] = dep_chan_data_5_0;
    assign token_in_vec_0[4] = token_5_0;
    assign in_chan_dep_vld_vec_0[5] = dep_chan_vld_7_0;
    assign in_chan_dep_data_vec_0[101 : 85] = dep_chan_data_7_0;
    assign token_in_vec_0[5] = token_7_0;
    assign in_chan_dep_vld_vec_0[6] = dep_chan_vld_16_0;
    assign in_chan_dep_data_vec_0[118 : 102] = dep_chan_data_16_0;
    assign token_in_vec_0[6] = token_16_0;
    assign dep_chan_vld_0_16 = out_chan_dep_vld_vec_0[0];
    assign dep_chan_data_0_16 = out_chan_dep_data_0;
    assign token_0_16 = token_out_vec_0[0];
    assign dep_chan_vld_0_5 = out_chan_dep_vld_vec_0[1];
    assign dep_chan_data_0_5 = out_chan_dep_data_0;
    assign token_0_5 = token_out_vec_0[1];
    assign dep_chan_vld_0_4 = out_chan_dep_vld_vec_0[2];
    assign dep_chan_data_0_4 = out_chan_dep_data_0;
    assign token_0_4 = token_out_vec_0[2];
    assign dep_chan_vld_0_1 = out_chan_dep_vld_vec_0[3];
    assign dep_chan_data_0_1 = out_chan_dep_data_0;
    assign token_0_1 = token_out_vec_0[3];
    assign dep_chan_vld_0_2 = out_chan_dep_vld_vec_0[4];
    assign dep_chan_data_0_2 = out_chan_dep_data_0;
    assign token_0_2 = token_out_vec_0[4];
    assign dep_chan_vld_0_3 = out_chan_dep_vld_vec_0[5];
    assign dep_chan_data_0_3 = out_chan_dep_data_0;
    assign token_0_3 = token_out_vec_0[5];
    assign dep_chan_vld_0_7 = out_chan_dep_vld_vec_0[6];
    assign dep_chan_data_0_7 = out_chan_dep_data_0;
    assign token_0_7 = token_out_vec_0[6];

    // Process: AESL_inst_top.Block_entry3_proc_U0
    AESL_deadlock_detect_unit #(17, 1, 9, 4) AESL_deadlock_detect_unit_1 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_1),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_1),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_1),
        .token_in_vec(token_in_vec_1),
        .dl_detect_in(dl_detect_out),
        .origin(origin[1]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_1),
        .out_chan_dep_data(out_chan_dep_data_1),
        .token_out_vec(token_out_vec_1),
        .dl_detect_out(dl_in_vec[1]));

    assign proc_1_data_FIFO_blk[0] = 1'b0;
    assign proc_1_data_PIPO_blk[0] = 1'b0;
    assign proc_1_start_FIFO_blk[0] = 1'b0;
    assign proc_1_TLF_FIFO_blk[0] = 1'b0;
    assign proc_1_input_sync_blk[0] = 1'b0 | (AESL_inst_top.ap_sync_Block_entry3_proc_U0_ap_ready & AESL_inst_top.Block_entry3_proc_U0.ap_idle & ~AESL_inst_top.ap_sync_entry_proc_U0_ap_ready);
    assign proc_1_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_1[0] = dl_detect_out ? proc_dep_vld_vec_1_reg[0] : (proc_1_data_FIFO_blk[0] | proc_1_data_PIPO_blk[0] | proc_1_start_FIFO_blk[0] | proc_1_TLF_FIFO_blk[0] | proc_1_input_sync_blk[0] | proc_1_output_sync_blk[0]);
    assign proc_1_data_FIFO_blk[1] = 1'b0;
    assign proc_1_data_PIPO_blk[1] = 1'b0;
    assign proc_1_start_FIFO_blk[1] = 1'b0;
    assign proc_1_TLF_FIFO_blk[1] = 1'b0;
    assign proc_1_input_sync_blk[1] = 1'b0 | (AESL_inst_top.ap_sync_Block_entry3_proc_U0_ap_ready & AESL_inst_top.Block_entry3_proc_U0.ap_idle & ~AESL_inst_top.ap_sync_ConvertBias_BN_U0_ap_ready);
    assign proc_1_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_1[1] = dl_detect_out ? proc_dep_vld_vec_1_reg[1] : (proc_1_data_FIFO_blk[1] | proc_1_data_PIPO_blk[1] | proc_1_start_FIFO_blk[1] | proc_1_TLF_FIFO_blk[1] | proc_1_input_sync_blk[1] | proc_1_output_sync_blk[1]);
    assign proc_1_data_FIFO_blk[2] = 1'b0;
    assign proc_1_data_PIPO_blk[2] = 1'b0;
    assign proc_1_start_FIFO_blk[2] = 1'b0;
    assign proc_1_TLF_FIFO_blk[2] = 1'b0;
    assign proc_1_input_sync_blk[2] = 1'b0 | (AESL_inst_top.ap_sync_Block_entry3_proc_U0_ap_ready & AESL_inst_top.Block_entry3_proc_U0.ap_idle & ~AESL_inst_top.ap_sync_ConvertInputToStream_U0_ap_ready);
    assign proc_1_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_1[2] = dl_detect_out ? proc_dep_vld_vec_1_reg[2] : (proc_1_data_FIFO_blk[2] | proc_1_data_PIPO_blk[2] | proc_1_start_FIFO_blk[2] | proc_1_TLF_FIFO_blk[2] | proc_1_input_sync_blk[2] | proc_1_output_sync_blk[2]);
    assign proc_1_data_FIFO_blk[3] = 1'b0;
    assign proc_1_data_PIPO_blk[3] = 1'b0;
    assign proc_1_start_FIFO_blk[3] = 1'b0;
    assign proc_1_TLF_FIFO_blk[3] = 1'b0;
    assign proc_1_input_sync_blk[3] = 1'b0 | (AESL_inst_top.ap_sync_Block_entry3_proc_U0_ap_ready & AESL_inst_top.Block_entry3_proc_U0.ap_idle & ~AESL_inst_top.ap_sync_ConvertWeightToStream_U0_ap_ready);
    assign proc_1_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_1[3] = dl_detect_out ? proc_dep_vld_vec_1_reg[3] : (proc_1_data_FIFO_blk[3] | proc_1_data_PIPO_blk[3] | proc_1_start_FIFO_blk[3] | proc_1_TLF_FIFO_blk[3] | proc_1_input_sync_blk[3] | proc_1_output_sync_blk[3]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_1_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_1_reg <= proc_dep_vld_vec_1;
        end
    end
    assign in_chan_dep_vld_vec_1[0] = dep_chan_vld_0_1;
    assign in_chan_dep_data_vec_1[16 : 0] = dep_chan_data_0_1;
    assign token_in_vec_1[0] = token_0_1;
    assign in_chan_dep_vld_vec_1[1] = dep_chan_vld_2_1;
    assign in_chan_dep_data_vec_1[33 : 17] = dep_chan_data_2_1;
    assign token_in_vec_1[1] = token_2_1;
    assign in_chan_dep_vld_vec_1[2] = dep_chan_vld_3_1;
    assign in_chan_dep_data_vec_1[50 : 34] = dep_chan_data_3_1;
    assign token_in_vec_1[2] = token_3_1;
    assign in_chan_dep_vld_vec_1[3] = dep_chan_vld_6_1;
    assign in_chan_dep_data_vec_1[67 : 51] = dep_chan_data_6_1;
    assign token_in_vec_1[3] = token_6_1;
    assign in_chan_dep_vld_vec_1[4] = dep_chan_vld_7_1;
    assign in_chan_dep_data_vec_1[84 : 68] = dep_chan_data_7_1;
    assign token_in_vec_1[4] = token_7_1;
    assign in_chan_dep_vld_vec_1[5] = dep_chan_vld_8_1;
    assign in_chan_dep_data_vec_1[101 : 85] = dep_chan_data_8_1;
    assign token_in_vec_1[5] = token_8_1;
    assign in_chan_dep_vld_vec_1[6] = dep_chan_vld_9_1;
    assign in_chan_dep_data_vec_1[118 : 102] = dep_chan_data_9_1;
    assign token_in_vec_1[6] = token_9_1;
    assign in_chan_dep_vld_vec_1[7] = dep_chan_vld_11_1;
    assign in_chan_dep_data_vec_1[135 : 119] = dep_chan_data_11_1;
    assign token_in_vec_1[7] = token_11_1;
    assign in_chan_dep_vld_vec_1[8] = dep_chan_vld_13_1;
    assign in_chan_dep_data_vec_1[152 : 136] = dep_chan_data_13_1;
    assign token_in_vec_1[8] = token_13_1;
    assign dep_chan_vld_1_0 = out_chan_dep_vld_vec_1[0];
    assign dep_chan_data_1_0 = out_chan_dep_data_1;
    assign token_1_0 = token_out_vec_1[0];
    assign dep_chan_vld_1_2 = out_chan_dep_vld_vec_1[1];
    assign dep_chan_data_1_2 = out_chan_dep_data_1;
    assign token_1_2 = token_out_vec_1[1];
    assign dep_chan_vld_1_3 = out_chan_dep_vld_vec_1[2];
    assign dep_chan_data_1_3 = out_chan_dep_data_1;
    assign token_1_3 = token_out_vec_1[2];
    assign dep_chan_vld_1_7 = out_chan_dep_vld_vec_1[3];
    assign dep_chan_data_1_7 = out_chan_dep_data_1;
    assign token_1_7 = token_out_vec_1[3];

    // Process: AESL_inst_top.ConvertBias_BN_U0
    AESL_deadlock_detect_unit #(17, 2, 6, 6) AESL_deadlock_detect_unit_2 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_2),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_2),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_2),
        .token_in_vec(token_in_vec_2),
        .dl_detect_in(dl_detect_out),
        .origin(origin[2]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_2),
        .out_chan_dep_data(out_chan_dep_data_2),
        .token_out_vec(token_out_vec_2),
        .dl_detect_out(dl_in_vec[2]));

    assign proc_2_data_FIFO_blk[0] = 1'b0 | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_0_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_1_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_2_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_3_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_4_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_5_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_6_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_7_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_8_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_9_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_10_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_11_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_12_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_13_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_14_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_15_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_16_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_17_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_18_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_19_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_20_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_21_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_22_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_23_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_24_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_25_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_26_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_27_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_28_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_29_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_30_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_31_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_32_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_33_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_34_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_35_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_36_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_37_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_38_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_39_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_40_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_41_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_42_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_43_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_44_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_45_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_46_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_47_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_48_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_49_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_50_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_51_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_52_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_53_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_54_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_55_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_56_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_57_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_58_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_59_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_60_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_61_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_62_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_63_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_64_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_65_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_66_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_67_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_68_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_69_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_70_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_71_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_72_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_73_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_74_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_75_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_76_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_77_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_78_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_79_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_80_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_81_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_82_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_83_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_84_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_85_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_86_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_87_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_88_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_89_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_90_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_91_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_92_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_93_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_94_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_95_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_96_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_97_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_98_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_99_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_100_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_101_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_102_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_103_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_104_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_105_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_106_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_107_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_108_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_109_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_110_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_111_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_112_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_113_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_114_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_115_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_116_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_117_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_118_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_119_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_120_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_121_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_122_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_123_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_124_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_125_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_126_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_127_blk_n);
    assign proc_2_data_PIPO_blk[0] = 1'b0;
    assign proc_2_start_FIFO_blk[0] = 1'b0 | (~AESL_inst_top.start_for_ConvBN_U0_U.if_full_n & AESL_inst_top.ConvertBias_BN_U0.ap_start & ~AESL_inst_top.ConvertBias_BN_U0.real_start & (trans_in_cnt_3 == trans_out_cnt_3) & ~AESL_inst_top.start_for_ConvBN_U0_U.if_read);
    assign proc_2_TLF_FIFO_blk[0] = 1'b0;
    assign proc_2_input_sync_blk[0] = 1'b0;
    assign proc_2_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_2[0] = dl_detect_out ? proc_dep_vld_vec_2_reg[0] : (proc_2_data_FIFO_blk[0] | proc_2_data_PIPO_blk[0] | proc_2_start_FIFO_blk[0] | proc_2_TLF_FIFO_blk[0] | proc_2_input_sync_blk[0] | proc_2_output_sync_blk[0]);
    assign proc_2_data_FIFO_blk[1] = 1'b0 | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_0_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_1_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_2_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_3_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_4_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_5_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_6_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_7_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_8_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_9_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_10_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_11_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_12_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_13_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_14_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_15_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_16_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_17_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_18_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_19_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_20_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_21_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_22_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_23_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_24_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_25_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_26_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_27_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_28_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_29_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_30_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_31_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_32_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_33_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_34_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_35_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_36_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_37_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_38_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_39_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_40_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_41_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_42_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_43_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_44_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_45_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_46_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_47_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_48_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_49_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_50_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_51_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_52_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_53_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_54_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_55_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_56_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_57_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_58_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_59_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_60_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_61_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_62_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_63_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_64_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_65_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_66_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_67_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_68_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_69_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_70_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_71_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_72_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_73_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_74_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_75_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_76_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_77_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_78_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_79_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_80_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_81_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_82_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_83_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_84_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_85_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_86_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_87_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_88_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_89_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_90_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_91_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_92_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_93_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_94_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_95_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_96_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_97_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_98_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_99_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_100_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_101_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_102_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_103_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_104_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_105_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_106_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_107_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_108_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_109_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_110_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_111_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_112_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_113_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_114_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_115_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_116_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_117_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_118_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_119_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_120_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_121_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_122_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_123_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_124_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_125_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_126_blk_n) | (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_127_blk_n);
    assign proc_2_data_PIPO_blk[1] = 1'b0;
    assign proc_2_start_FIFO_blk[1] = 1'b0 | (~AESL_inst_top.start_for_ConvBias_U0_U.if_full_n & AESL_inst_top.ConvertBias_BN_U0.ap_start & ~AESL_inst_top.ConvertBias_BN_U0.real_start & (trans_in_cnt_3 == trans_out_cnt_3) & ~AESL_inst_top.start_for_ConvBias_U0_U.if_read);
    assign proc_2_TLF_FIFO_blk[1] = 1'b0;
    assign proc_2_input_sync_blk[1] = 1'b0;
    assign proc_2_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_2[1] = dl_detect_out ? proc_dep_vld_vec_2_reg[1] : (proc_2_data_FIFO_blk[1] | proc_2_data_PIPO_blk[1] | proc_2_start_FIFO_blk[1] | proc_2_TLF_FIFO_blk[1] | proc_2_input_sync_blk[1] | proc_2_output_sync_blk[1]);
    assign proc_2_data_FIFO_blk[2] = 1'b0;
    assign proc_2_data_PIPO_blk[2] = 1'b0;
    assign proc_2_start_FIFO_blk[2] = 1'b0;
    assign proc_2_TLF_FIFO_blk[2] = 1'b0;
    assign proc_2_input_sync_blk[2] = 1'b0 | (AESL_inst_top.ap_sync_ConvertBias_BN_U0_ap_ready & AESL_inst_top.ConvertBias_BN_U0.ap_idle & ~AESL_inst_top.ap_sync_entry_proc_U0_ap_ready);
    assign proc_2_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_2[2] = dl_detect_out ? proc_dep_vld_vec_2_reg[2] : (proc_2_data_FIFO_blk[2] | proc_2_data_PIPO_blk[2] | proc_2_start_FIFO_blk[2] | proc_2_TLF_FIFO_blk[2] | proc_2_input_sync_blk[2] | proc_2_output_sync_blk[2]);
    assign proc_2_data_FIFO_blk[3] = 1'b0;
    assign proc_2_data_PIPO_blk[3] = 1'b0;
    assign proc_2_start_FIFO_blk[3] = 1'b0;
    assign proc_2_TLF_FIFO_blk[3] = 1'b0;
    assign proc_2_input_sync_blk[3] = 1'b0 | (AESL_inst_top.ap_sync_ConvertBias_BN_U0_ap_ready & AESL_inst_top.ConvertBias_BN_U0.ap_idle & ~AESL_inst_top.ap_sync_Block_entry3_proc_U0_ap_ready);
    assign proc_2_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_2[3] = dl_detect_out ? proc_dep_vld_vec_2_reg[3] : (proc_2_data_FIFO_blk[3] | proc_2_data_PIPO_blk[3] | proc_2_start_FIFO_blk[3] | proc_2_TLF_FIFO_blk[3] | proc_2_input_sync_blk[3] | proc_2_output_sync_blk[3]);
    assign proc_2_data_FIFO_blk[4] = 1'b0;
    assign proc_2_data_PIPO_blk[4] = 1'b0;
    assign proc_2_start_FIFO_blk[4] = 1'b0;
    assign proc_2_TLF_FIFO_blk[4] = 1'b0;
    assign proc_2_input_sync_blk[4] = 1'b0 | (AESL_inst_top.ap_sync_ConvertBias_BN_U0_ap_ready & AESL_inst_top.ConvertBias_BN_U0.ap_idle & ~AESL_inst_top.ap_sync_ConvertInputToStream_U0_ap_ready);
    assign proc_2_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_2[4] = dl_detect_out ? proc_dep_vld_vec_2_reg[4] : (proc_2_data_FIFO_blk[4] | proc_2_data_PIPO_blk[4] | proc_2_start_FIFO_blk[4] | proc_2_TLF_FIFO_blk[4] | proc_2_input_sync_blk[4] | proc_2_output_sync_blk[4]);
    assign proc_2_data_FIFO_blk[5] = 1'b0;
    assign proc_2_data_PIPO_blk[5] = 1'b0;
    assign proc_2_start_FIFO_blk[5] = 1'b0;
    assign proc_2_TLF_FIFO_blk[5] = 1'b0;
    assign proc_2_input_sync_blk[5] = 1'b0 | (AESL_inst_top.ap_sync_ConvertBias_BN_U0_ap_ready & AESL_inst_top.ConvertBias_BN_U0.ap_idle & ~AESL_inst_top.ap_sync_ConvertWeightToStream_U0_ap_ready);
    assign proc_2_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_2[5] = dl_detect_out ? proc_dep_vld_vec_2_reg[5] : (proc_2_data_FIFO_blk[5] | proc_2_data_PIPO_blk[5] | proc_2_start_FIFO_blk[5] | proc_2_TLF_FIFO_blk[5] | proc_2_input_sync_blk[5] | proc_2_output_sync_blk[5]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_2_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_2_reg <= proc_dep_vld_vec_2;
        end
    end
    assign in_chan_dep_vld_vec_2[0] = dep_chan_vld_0_2;
    assign in_chan_dep_data_vec_2[16 : 0] = dep_chan_data_0_2;
    assign token_in_vec_2[0] = token_0_2;
    assign in_chan_dep_vld_vec_2[1] = dep_chan_vld_1_2;
    assign in_chan_dep_data_vec_2[33 : 17] = dep_chan_data_1_2;
    assign token_in_vec_2[1] = token_1_2;
    assign in_chan_dep_vld_vec_2[2] = dep_chan_vld_3_2;
    assign in_chan_dep_data_vec_2[50 : 34] = dep_chan_data_3_2;
    assign token_in_vec_2[2] = token_3_2;
    assign in_chan_dep_vld_vec_2[3] = dep_chan_vld_7_2;
    assign in_chan_dep_data_vec_2[67 : 51] = dep_chan_data_7_2;
    assign token_in_vec_2[3] = token_7_2;
    assign in_chan_dep_vld_vec_2[4] = dep_chan_vld_14_2;
    assign in_chan_dep_data_vec_2[84 : 68] = dep_chan_data_14_2;
    assign token_in_vec_2[4] = token_14_2;
    assign in_chan_dep_vld_vec_2[5] = dep_chan_vld_15_2;
    assign in_chan_dep_data_vec_2[101 : 85] = dep_chan_data_15_2;
    assign token_in_vec_2[5] = token_15_2;
    assign dep_chan_vld_2_15 = out_chan_dep_vld_vec_2[0];
    assign dep_chan_data_2_15 = out_chan_dep_data_2;
    assign token_2_15 = token_out_vec_2[0];
    assign dep_chan_vld_2_14 = out_chan_dep_vld_vec_2[1];
    assign dep_chan_data_2_14 = out_chan_dep_data_2;
    assign token_2_14 = token_out_vec_2[1];
    assign dep_chan_vld_2_0 = out_chan_dep_vld_vec_2[2];
    assign dep_chan_data_2_0 = out_chan_dep_data_2;
    assign token_2_0 = token_out_vec_2[2];
    assign dep_chan_vld_2_1 = out_chan_dep_vld_vec_2[3];
    assign dep_chan_data_2_1 = out_chan_dep_data_2;
    assign token_2_1 = token_out_vec_2[3];
    assign dep_chan_vld_2_3 = out_chan_dep_vld_vec_2[4];
    assign dep_chan_data_2_3 = out_chan_dep_data_2;
    assign token_2_3 = token_out_vec_2[4];
    assign dep_chan_vld_2_7 = out_chan_dep_vld_vec_2[5];
    assign dep_chan_data_2_7 = out_chan_dep_data_2;
    assign token_2_7 = token_out_vec_2[5];

    // Process: AESL_inst_top.ConvertInputToStream_U0
    AESL_deadlock_detect_unit #(17, 3, 6, 6) AESL_deadlock_detect_unit_3 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_3),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_3),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_3),
        .token_in_vec(token_in_vec_3),
        .dl_detect_in(dl_detect_out),
        .origin(origin[3]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_3),
        .out_chan_dep_data(out_chan_dep_data_3),
        .token_out_vec(token_out_vec_3),
        .dl_detect_out(dl_in_vec[3]));

    assign proc_3_data_FIFO_blk[0] = 1'b0 | (~AESL_inst_top.ConvertInputToStream_U0.grp_ConvertInputToStream_Pipeline_VITIS_LOOP_19_1_VITIS_LOOP_22_2_VITIS_LOOP_25_3_VI_fu_166.conv_a_blk_n) | (~AESL_inst_top.ConvertInputToStream_U0.R_c46_blk_n) | (~AESL_inst_top.ConvertInputToStream_U0.C_c48_blk_n) | (~AESL_inst_top.ConvertInputToStream_U0.N_c51_blk_n) | (~AESL_inst_top.ConvertInputToStream_U0.M_c56_blk_n) | (~AESL_inst_top.ConvertInputToStream_U0.mode_c72_blk_n);
    assign proc_3_data_PIPO_blk[0] = 1'b0;
    assign proc_3_start_FIFO_blk[0] = 1'b0;
    assign proc_3_TLF_FIFO_blk[0] = 1'b0;
    assign proc_3_input_sync_blk[0] = 1'b0;
    assign proc_3_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_3[0] = dl_detect_out ? proc_dep_vld_vec_3_reg[0] : (proc_3_data_FIFO_blk[0] | proc_3_data_PIPO_blk[0] | proc_3_start_FIFO_blk[0] | proc_3_TLF_FIFO_blk[0] | proc_3_input_sync_blk[0] | proc_3_output_sync_blk[0]);
    assign proc_3_data_FIFO_blk[1] = 1'b0 | (~AESL_inst_top.ConvertInputToStream_U0.grp_ConvertInputToStream_Pipeline_VITIS_LOOP_40_5_VITIS_LOOP_43_6_VITIS_LOOP_46_7_fu_154.mm_a_blk_n);
    assign proc_3_data_PIPO_blk[1] = 1'b0;
    assign proc_3_start_FIFO_blk[1] = 1'b0;
    assign proc_3_TLF_FIFO_blk[1] = 1'b0;
    assign proc_3_input_sync_blk[1] = 1'b0;
    assign proc_3_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_3[1] = dl_detect_out ? proc_dep_vld_vec_3_reg[1] : (proc_3_data_FIFO_blk[1] | proc_3_data_PIPO_blk[1] | proc_3_start_FIFO_blk[1] | proc_3_TLF_FIFO_blk[1] | proc_3_input_sync_blk[1] | proc_3_output_sync_blk[1]);
    assign proc_3_data_FIFO_blk[2] = 1'b0;
    assign proc_3_data_PIPO_blk[2] = 1'b0;
    assign proc_3_start_FIFO_blk[2] = 1'b0;
    assign proc_3_TLF_FIFO_blk[2] = 1'b0;
    assign proc_3_input_sync_blk[2] = 1'b0 | (AESL_inst_top.ap_sync_ConvertInputToStream_U0_ap_ready & AESL_inst_top.ConvertInputToStream_U0.ap_idle & ~AESL_inst_top.ap_sync_entry_proc_U0_ap_ready);
    assign proc_3_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_3[2] = dl_detect_out ? proc_dep_vld_vec_3_reg[2] : (proc_3_data_FIFO_blk[2] | proc_3_data_PIPO_blk[2] | proc_3_start_FIFO_blk[2] | proc_3_TLF_FIFO_blk[2] | proc_3_input_sync_blk[2] | proc_3_output_sync_blk[2]);
    assign proc_3_data_FIFO_blk[3] = 1'b0;
    assign proc_3_data_PIPO_blk[3] = 1'b0;
    assign proc_3_start_FIFO_blk[3] = 1'b0;
    assign proc_3_TLF_FIFO_blk[3] = 1'b0;
    assign proc_3_input_sync_blk[3] = 1'b0 | (AESL_inst_top.ap_sync_ConvertInputToStream_U0_ap_ready & AESL_inst_top.ConvertInputToStream_U0.ap_idle & ~AESL_inst_top.ap_sync_Block_entry3_proc_U0_ap_ready);
    assign proc_3_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_3[3] = dl_detect_out ? proc_dep_vld_vec_3_reg[3] : (proc_3_data_FIFO_blk[3] | proc_3_data_PIPO_blk[3] | proc_3_start_FIFO_blk[3] | proc_3_TLF_FIFO_blk[3] | proc_3_input_sync_blk[3] | proc_3_output_sync_blk[3]);
    assign proc_3_data_FIFO_blk[4] = 1'b0;
    assign proc_3_data_PIPO_blk[4] = 1'b0;
    assign proc_3_start_FIFO_blk[4] = 1'b0;
    assign proc_3_TLF_FIFO_blk[4] = 1'b0;
    assign proc_3_input_sync_blk[4] = 1'b0 | (AESL_inst_top.ap_sync_ConvertInputToStream_U0_ap_ready & AESL_inst_top.ConvertInputToStream_U0.ap_idle & ~AESL_inst_top.ap_sync_ConvertBias_BN_U0_ap_ready);
    assign proc_3_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_3[4] = dl_detect_out ? proc_dep_vld_vec_3_reg[4] : (proc_3_data_FIFO_blk[4] | proc_3_data_PIPO_blk[4] | proc_3_start_FIFO_blk[4] | proc_3_TLF_FIFO_blk[4] | proc_3_input_sync_blk[4] | proc_3_output_sync_blk[4]);
    assign proc_3_data_FIFO_blk[5] = 1'b0;
    assign proc_3_data_PIPO_blk[5] = 1'b0;
    assign proc_3_start_FIFO_blk[5] = 1'b0;
    assign proc_3_TLF_FIFO_blk[5] = 1'b0;
    assign proc_3_input_sync_blk[5] = 1'b0 | (AESL_inst_top.ap_sync_ConvertInputToStream_U0_ap_ready & AESL_inst_top.ConvertInputToStream_U0.ap_idle & ~AESL_inst_top.ap_sync_ConvertWeightToStream_U0_ap_ready);
    assign proc_3_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_3[5] = dl_detect_out ? proc_dep_vld_vec_3_reg[5] : (proc_3_data_FIFO_blk[5] | proc_3_data_PIPO_blk[5] | proc_3_start_FIFO_blk[5] | proc_3_TLF_FIFO_blk[5] | proc_3_input_sync_blk[5] | proc_3_output_sync_blk[5]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_3_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_3_reg <= proc_dep_vld_vec_3;
        end
    end
    assign in_chan_dep_vld_vec_3[0] = dep_chan_vld_0_3;
    assign in_chan_dep_data_vec_3[16 : 0] = dep_chan_data_0_3;
    assign token_in_vec_3[0] = token_0_3;
    assign in_chan_dep_vld_vec_3[1] = dep_chan_vld_1_3;
    assign in_chan_dep_data_vec_3[33 : 17] = dep_chan_data_1_3;
    assign token_in_vec_3[1] = token_1_3;
    assign in_chan_dep_vld_vec_3[2] = dep_chan_vld_2_3;
    assign in_chan_dep_data_vec_3[50 : 34] = dep_chan_data_2_3;
    assign token_in_vec_3[2] = token_2_3;
    assign in_chan_dep_vld_vec_3[3] = dep_chan_vld_4_3;
    assign in_chan_dep_data_vec_3[67 : 51] = dep_chan_data_4_3;
    assign token_in_vec_3[3] = token_4_3;
    assign in_chan_dep_vld_vec_3[4] = dep_chan_vld_6_3;
    assign in_chan_dep_data_vec_3[84 : 68] = dep_chan_data_6_3;
    assign token_in_vec_3[4] = token_6_3;
    assign in_chan_dep_vld_vec_3[5] = dep_chan_vld_7_3;
    assign in_chan_dep_data_vec_3[101 : 85] = dep_chan_data_7_3;
    assign token_in_vec_3[5] = token_7_3;
    assign dep_chan_vld_3_4 = out_chan_dep_vld_vec_3[0];
    assign dep_chan_data_3_4 = out_chan_dep_data_3;
    assign token_3_4 = token_out_vec_3[0];
    assign dep_chan_vld_3_6 = out_chan_dep_vld_vec_3[1];
    assign dep_chan_data_3_6 = out_chan_dep_data_3;
    assign token_3_6 = token_out_vec_3[1];
    assign dep_chan_vld_3_0 = out_chan_dep_vld_vec_3[2];
    assign dep_chan_data_3_0 = out_chan_dep_data_3;
    assign token_3_0 = token_out_vec_3[2];
    assign dep_chan_vld_3_1 = out_chan_dep_vld_vec_3[3];
    assign dep_chan_data_3_1 = out_chan_dep_data_3;
    assign token_3_1 = token_out_vec_3[3];
    assign dep_chan_vld_3_2 = out_chan_dep_vld_vec_3[4];
    assign dep_chan_data_3_2 = out_chan_dep_data_3;
    assign token_3_2 = token_out_vec_3[4];
    assign dep_chan_vld_3_7 = out_chan_dep_vld_vec_3[5];
    assign dep_chan_data_3_7 = out_chan_dep_data_3;
    assign token_3_7 = token_out_vec_3[5];

    // Process: AESL_inst_top.Padding_U0
    AESL_deadlock_detect_unit #(17, 4, 3, 3) AESL_deadlock_detect_unit_4 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_4),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_4),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_4),
        .token_in_vec(token_in_vec_4),
        .dl_detect_in(dl_detect_out),
        .origin(origin[4]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_4),
        .out_chan_dep_data(out_chan_dep_data_4),
        .token_out_vec(token_out_vec_4),
        .dl_detect_out(dl_in_vec[4]));

    assign proc_4_data_FIFO_blk[0] = 1'b0 | (~AESL_inst_top.Padding_U0.grp_Padding_Pipeline_VITIS_LOOP_62_1_VITIS_LOOP_65_2_VITIS_LOOP_68_3_VITIS_LOOP_71_4_fu_152.conv_a_blk_n) | (~AESL_inst_top.Padding_U0.R_blk_n) | (~AESL_inst_top.Padding_U0.C_blk_n) | (~AESL_inst_top.Padding_U0.N_blk_n) | (~AESL_inst_top.Padding_U0.M_blk_n) | (~AESL_inst_top.Padding_U0.mode_blk_n);
    assign proc_4_data_PIPO_blk[0] = 1'b0;
    assign proc_4_start_FIFO_blk[0] = 1'b0;
    assign proc_4_TLF_FIFO_blk[0] = 1'b0;
    assign proc_4_input_sync_blk[0] = 1'b0;
    assign proc_4_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_4[0] = dl_detect_out ? proc_dep_vld_vec_4_reg[0] : (proc_4_data_FIFO_blk[0] | proc_4_data_PIPO_blk[0] | proc_4_start_FIFO_blk[0] | proc_4_TLF_FIFO_blk[0] | proc_4_input_sync_blk[0] | proc_4_output_sync_blk[0]);
    assign proc_4_data_FIFO_blk[1] = 1'b0 | (~AESL_inst_top.Padding_U0.grp_Padding_Pipeline_VITIS_LOOP_62_1_VITIS_LOOP_65_2_VITIS_LOOP_68_3_VITIS_LOOP_71_4_fu_152.conv3_samepad_blk_n) | (~AESL_inst_top.Padding_U0.R_c45_blk_n) | (~AESL_inst_top.Padding_U0.C_c47_blk_n) | (~AESL_inst_top.Padding_U0.N_c50_blk_n) | (~AESL_inst_top.Padding_U0.M_c55_blk_n) | (~AESL_inst_top.Padding_U0.P_c59_blk_n) | (~AESL_inst_top.Padding_U0.mode_c71_blk_n);
    assign proc_4_data_PIPO_blk[1] = 1'b0;
    assign proc_4_start_FIFO_blk[1] = 1'b0;
    assign proc_4_TLF_FIFO_blk[1] = 1'b0;
    assign proc_4_input_sync_blk[1] = 1'b0;
    assign proc_4_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_4[1] = dl_detect_out ? proc_dep_vld_vec_4_reg[1] : (proc_4_data_FIFO_blk[1] | proc_4_data_PIPO_blk[1] | proc_4_start_FIFO_blk[1] | proc_4_TLF_FIFO_blk[1] | proc_4_input_sync_blk[1] | proc_4_output_sync_blk[1]);
    assign proc_4_data_FIFO_blk[2] = 1'b0 | (~AESL_inst_top.Padding_U0.P_blk_n);
    assign proc_4_data_PIPO_blk[2] = 1'b0;
    assign proc_4_start_FIFO_blk[2] = 1'b0 | (~AESL_inst_top.start_for_Padding_U0_U.if_empty_n & AESL_inst_top.Padding_U0.ap_idle & ~AESL_inst_top.start_for_Padding_U0_U.if_write);
    assign proc_4_TLF_FIFO_blk[2] = 1'b0;
    assign proc_4_input_sync_blk[2] = 1'b0;
    assign proc_4_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_4[2] = dl_detect_out ? proc_dep_vld_vec_4_reg[2] : (proc_4_data_FIFO_blk[2] | proc_4_data_PIPO_blk[2] | proc_4_start_FIFO_blk[2] | proc_4_TLF_FIFO_blk[2] | proc_4_input_sync_blk[2] | proc_4_output_sync_blk[2]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_4_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_4_reg <= proc_dep_vld_vec_4;
        end
    end
    assign in_chan_dep_vld_vec_4[0] = dep_chan_vld_0_4;
    assign in_chan_dep_data_vec_4[16 : 0] = dep_chan_data_0_4;
    assign token_in_vec_4[0] = token_0_4;
    assign in_chan_dep_vld_vec_4[1] = dep_chan_vld_3_4;
    assign in_chan_dep_data_vec_4[33 : 17] = dep_chan_data_3_4;
    assign token_in_vec_4[1] = token_3_4;
    assign in_chan_dep_vld_vec_4[2] = dep_chan_vld_5_4;
    assign in_chan_dep_data_vec_4[50 : 34] = dep_chan_data_5_4;
    assign token_in_vec_4[2] = token_5_4;
    assign dep_chan_vld_4_3 = out_chan_dep_vld_vec_4[0];
    assign dep_chan_data_4_3 = out_chan_dep_data_4;
    assign token_4_3 = token_out_vec_4[0];
    assign dep_chan_vld_4_5 = out_chan_dep_vld_vec_4[1];
    assign dep_chan_data_4_5 = out_chan_dep_data_4;
    assign token_4_5 = token_out_vec_4[1];
    assign dep_chan_vld_4_0 = out_chan_dep_vld_vec_4[2];
    assign dep_chan_data_4_0 = out_chan_dep_data_4;
    assign token_4_0 = token_out_vec_4[2];

    // Process: AESL_inst_top.Sliding_U0
    AESL_deadlock_detect_unit #(17, 5, 6, 6) AESL_deadlock_detect_unit_5 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_5),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_5),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_5),
        .token_in_vec(token_in_vec_5),
        .dl_detect_in(dl_detect_out),
        .origin(origin[5]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_5),
        .out_chan_dep_data(out_chan_dep_data_5),
        .token_out_vec(token_out_vec_5),
        .dl_detect_out(dl_in_vec[5]));

    assign proc_5_data_FIFO_blk[0] = 1'b0 | (~AESL_inst_top.Sliding_U0.grp_Sliding_Pipeline_VITIS_LOOP_114_1_VITIS_LOOP_117_2_fu_192.conv3_samepad_blk_n) | (~AESL_inst_top.Sliding_U0.R_blk_n) | (~AESL_inst_top.Sliding_U0.C_blk_n) | (~AESL_inst_top.Sliding_U0.N_blk_n) | (~AESL_inst_top.Sliding_U0.M_blk_n) | (~AESL_inst_top.Sliding_U0.P_blk_n) | (~AESL_inst_top.Sliding_U0.mode_blk_n);
    assign proc_5_data_PIPO_blk[0] = 1'b0;
    assign proc_5_start_FIFO_blk[0] = 1'b0;
    assign proc_5_TLF_FIFO_blk[0] = 1'b0;
    assign proc_5_input_sync_blk[0] = 1'b0;
    assign proc_5_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_5[0] = dl_detect_out ? proc_dep_vld_vec_5_reg[0] : (proc_5_data_FIFO_blk[0] | proc_5_data_PIPO_blk[0] | proc_5_start_FIFO_blk[0] | proc_5_TLF_FIFO_blk[0] | proc_5_input_sync_blk[0] | proc_5_output_sync_blk[0]);
    assign proc_5_data_FIFO_blk[1] = 1'b0 | (~AESL_inst_top.Sliding_U0.grp_Sliding_Pipeline_VITIS_LOOP_114_1_VITIS_LOOP_117_2_fu_192.conv3_sild_blk_n) | (~AESL_inst_top.Sliding_U0.mode_c70_blk_n);
    assign proc_5_data_PIPO_blk[1] = 1'b0;
    assign proc_5_start_FIFO_blk[1] = 1'b0;
    assign proc_5_TLF_FIFO_blk[1] = 1'b0;
    assign proc_5_input_sync_blk[1] = 1'b0;
    assign proc_5_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_5[1] = dl_detect_out ? proc_dep_vld_vec_5_reg[1] : (proc_5_data_FIFO_blk[1] | proc_5_data_PIPO_blk[1] | proc_5_start_FIFO_blk[1] | proc_5_TLF_FIFO_blk[1] | proc_5_input_sync_blk[1] | proc_5_output_sync_blk[1]);
    assign proc_5_data_FIFO_blk[2] = 1'b0 | (~AESL_inst_top.Sliding_U0.K_blk_n) | (~AESL_inst_top.Sliding_U0.S_blk_n);
    assign proc_5_data_PIPO_blk[2] = 1'b0;
    assign proc_5_start_FIFO_blk[2] = 1'b0 | (~AESL_inst_top.start_for_Sliding_U0_U.if_empty_n & AESL_inst_top.Sliding_U0.ap_idle & ~AESL_inst_top.start_for_Sliding_U0_U.if_write);
    assign proc_5_TLF_FIFO_blk[2] = 1'b0;
    assign proc_5_input_sync_blk[2] = 1'b0;
    assign proc_5_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_5[2] = dl_detect_out ? proc_dep_vld_vec_5_reg[2] : (proc_5_data_FIFO_blk[2] | proc_5_data_PIPO_blk[2] | proc_5_start_FIFO_blk[2] | proc_5_TLF_FIFO_blk[2] | proc_5_input_sync_blk[2] | proc_5_output_sync_blk[2]);
    assign proc_5_data_FIFO_blk[3] = 1'b0 | (~AESL_inst_top.Sliding_U0.R_c44_blk_n) | (~AESL_inst_top.Sliding_U0.N_c49_blk_n);
    assign proc_5_data_PIPO_blk[3] = 1'b0;
    assign proc_5_start_FIFO_blk[3] = 1'b0 | (~AESL_inst_top.start_for_ConvertToOutStream_U0_U.if_full_n & AESL_inst_top.Sliding_U0.ap_start & ~AESL_inst_top.Sliding_U0.real_start & (trans_in_cnt_2 == trans_out_cnt_2) & ~AESL_inst_top.start_for_ConvertToOutStream_U0_U.if_read);
    assign proc_5_TLF_FIFO_blk[3] = 1'b0;
    assign proc_5_input_sync_blk[3] = 1'b0;
    assign proc_5_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_5[3] = dl_detect_out ? proc_dep_vld_vec_5_reg[3] : (proc_5_data_FIFO_blk[3] | proc_5_data_PIPO_blk[3] | proc_5_start_FIFO_blk[3] | proc_5_TLF_FIFO_blk[3] | proc_5_input_sync_blk[3] | proc_5_output_sync_blk[3]);
    assign proc_5_data_FIFO_blk[4] = 1'b0 | (~AESL_inst_top.Sliding_U0.C_c_blk_n) | (~AESL_inst_top.Sliding_U0.P_c_blk_n) | (~AESL_inst_top.Sliding_U0.S_c_blk_n);
    assign proc_5_data_PIPO_blk[4] = 1'b0;
    assign proc_5_start_FIFO_blk[4] = 1'b0;
    assign proc_5_TLF_FIFO_blk[4] = 1'b0;
    assign proc_5_input_sync_blk[4] = 1'b0;
    assign proc_5_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_5[4] = dl_detect_out ? proc_dep_vld_vec_5_reg[4] : (proc_5_data_FIFO_blk[4] | proc_5_data_PIPO_blk[4] | proc_5_start_FIFO_blk[4] | proc_5_TLF_FIFO_blk[4] | proc_5_input_sync_blk[4] | proc_5_output_sync_blk[4]);
    assign proc_5_data_FIFO_blk[5] = 1'b0 | (~AESL_inst_top.Sliding_U0.M_c54_blk_n) | (~AESL_inst_top.Sliding_U0.K_c57_blk_n);
    assign proc_5_data_PIPO_blk[5] = 1'b0;
    assign proc_5_start_FIFO_blk[5] = 1'b0;
    assign proc_5_TLF_FIFO_blk[5] = 1'b0;
    assign proc_5_input_sync_blk[5] = 1'b0;
    assign proc_5_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_5[5] = dl_detect_out ? proc_dep_vld_vec_5_reg[5] : (proc_5_data_FIFO_blk[5] | proc_5_data_PIPO_blk[5] | proc_5_start_FIFO_blk[5] | proc_5_TLF_FIFO_blk[5] | proc_5_input_sync_blk[5] | proc_5_output_sync_blk[5]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_5_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_5_reg <= proc_dep_vld_vec_5;
        end
    end
    assign in_chan_dep_vld_vec_5[0] = dep_chan_vld_0_5;
    assign in_chan_dep_data_vec_5[16 : 0] = dep_chan_data_0_5;
    assign token_in_vec_5[0] = token_0_5;
    assign in_chan_dep_vld_vec_5[1] = dep_chan_vld_4_5;
    assign in_chan_dep_data_vec_5[33 : 17] = dep_chan_data_4_5;
    assign token_in_vec_5[1] = token_4_5;
    assign in_chan_dep_vld_vec_5[2] = dep_chan_vld_6_5;
    assign in_chan_dep_data_vec_5[50 : 34] = dep_chan_data_6_5;
    assign token_in_vec_5[2] = token_6_5;
    assign in_chan_dep_vld_vec_5[3] = dep_chan_vld_12_5;
    assign in_chan_dep_data_vec_5[67 : 51] = dep_chan_data_12_5;
    assign token_in_vec_5[3] = token_12_5;
    assign in_chan_dep_vld_vec_5[4] = dep_chan_vld_13_5;
    assign in_chan_dep_data_vec_5[84 : 68] = dep_chan_data_13_5;
    assign token_in_vec_5[4] = token_13_5;
    assign in_chan_dep_vld_vec_5[5] = dep_chan_vld_16_5;
    assign in_chan_dep_data_vec_5[101 : 85] = dep_chan_data_16_5;
    assign token_in_vec_5[5] = token_16_5;
    assign dep_chan_vld_5_4 = out_chan_dep_vld_vec_5[0];
    assign dep_chan_data_5_4 = out_chan_dep_data_5;
    assign token_5_4 = token_out_vec_5[0];
    assign dep_chan_vld_5_6 = out_chan_dep_vld_vec_5[1];
    assign dep_chan_data_5_6 = out_chan_dep_data_5;
    assign token_5_6 = token_out_vec_5[1];
    assign dep_chan_vld_5_0 = out_chan_dep_vld_vec_5[2];
    assign dep_chan_data_5_0 = out_chan_dep_data_5;
    assign token_5_0 = token_out_vec_5[2];
    assign dep_chan_vld_5_12 = out_chan_dep_vld_vec_5[3];
    assign dep_chan_data_5_12 = out_chan_dep_data_5;
    assign token_5_12 = token_out_vec_5[3];
    assign dep_chan_vld_5_16 = out_chan_dep_vld_vec_5[4];
    assign dep_chan_data_5_16 = out_chan_dep_data_5;
    assign token_5_16 = token_out_vec_5[4];
    assign dep_chan_vld_5_13 = out_chan_dep_vld_vec_5[5];
    assign dep_chan_data_5_13 = out_chan_dep_data_5;
    assign token_5_13 = token_out_vec_5[5];

    // Process: AESL_inst_top.ConvertInputToArray_U0
    AESL_deadlock_detect_unit #(17, 6, 3, 4) AESL_deadlock_detect_unit_6 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_6),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_6),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_6),
        .token_in_vec(token_in_vec_6),
        .dl_detect_in(dl_detect_out),
        .origin(origin[6]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_6),
        .out_chan_dep_data(out_chan_dep_data_6),
        .token_out_vec(token_out_vec_6),
        .dl_detect_out(dl_in_vec[6]));

    assign proc_6_data_FIFO_blk[0] = 1'b0 | (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.conv3_sild_blk_n) | (~AESL_inst_top.ConvertInputToArray_U0.mode_blk_n);
    assign proc_6_data_PIPO_blk[0] = 1'b0;
    assign proc_6_start_FIFO_blk[0] = 1'b0;
    assign proc_6_TLF_FIFO_blk[0] = 1'b0;
    assign proc_6_input_sync_blk[0] = 1'b0;
    assign proc_6_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_6[0] = dl_detect_out ? proc_dep_vld_vec_6_reg[0] : (proc_6_data_FIFO_blk[0] | proc_6_data_PIPO_blk[0] | proc_6_start_FIFO_blk[0] | proc_6_TLF_FIFO_blk[0] | proc_6_input_sync_blk[0] | proc_6_output_sync_blk[0]);
    assign proc_6_data_FIFO_blk[1] = 1'b0 | (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.mm_a_blk_n);
    assign proc_6_data_PIPO_blk[1] = 1'b0;
    assign proc_6_start_FIFO_blk[1] = 1'b0;
    assign proc_6_TLF_FIFO_blk[1] = 1'b0;
    assign proc_6_input_sync_blk[1] = 1'b0;
    assign proc_6_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_6[1] = dl_detect_out ? proc_dep_vld_vec_6_reg[1] : (proc_6_data_FIFO_blk[1] | proc_6_data_PIPO_blk[1] | proc_6_start_FIFO_blk[1] | proc_6_TLF_FIFO_blk[1] | proc_6_input_sync_blk[1] | proc_6_output_sync_blk[1]);
    assign proc_6_data_FIFO_blk[2] = 1'b0 | (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.fifo_SA_A_blk_n) | (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.fifo_SA_A_1_blk_n) | (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.fifo_SA_A_2_blk_n) | (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.fifo_SA_A_3_blk_n) | (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.fifo_SA_A_4_blk_n) | (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.fifo_SA_A_5_blk_n) | (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.fifo_SA_A_6_blk_n) | (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.fifo_SA_A_7_blk_n) | (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.fifo_SA_A_8_blk_n) | (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.fifo_SA_A_9_blk_n) | (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.fifo_SA_A_10_blk_n) | (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.fifo_SA_A_11_blk_n) | (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.fifo_SA_A_12_blk_n) | (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.fifo_SA_A_13_blk_n) | (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.fifo_SA_A_14_blk_n) | (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.fifo_SA_A_15_blk_n) | (~AESL_inst_top.ConvertInputToArray_U0.num_a_sa_2_loc_c42_blk_n) | (~AESL_inst_top.ConvertInputToArray_U0.mode_c66_blk_n);
    assign proc_6_data_PIPO_blk[2] = 1'b0;
    assign proc_6_start_FIFO_blk[2] = 1'b0;
    assign proc_6_TLF_FIFO_blk[2] = 1'b0;
    assign proc_6_input_sync_blk[2] = 1'b0;
    assign proc_6_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_6[2] = dl_detect_out ? proc_dep_vld_vec_6_reg[2] : (proc_6_data_FIFO_blk[2] | proc_6_data_PIPO_blk[2] | proc_6_start_FIFO_blk[2] | proc_6_TLF_FIFO_blk[2] | proc_6_input_sync_blk[2] | proc_6_output_sync_blk[2]);
    assign proc_6_data_FIFO_blk[3] = 1'b0;
    assign proc_6_data_PIPO_blk[3] = 1'b0;
    assign proc_6_start_FIFO_blk[3] = 1'b0;
    assign proc_6_TLF_FIFO_blk[3] = 1'b0 | (~AESL_inst_top.num_a_sa_2_loc_c43_channel_U.if_empty_n & AESL_inst_top.ConvertInputToArray_U0.ap_idle & ~AESL_inst_top.num_a_sa_2_loc_c43_channel_U.if_write);
    assign proc_6_input_sync_blk[3] = 1'b0;
    assign proc_6_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_6[3] = dl_detect_out ? proc_dep_vld_vec_6_reg[3] : (proc_6_data_FIFO_blk[3] | proc_6_data_PIPO_blk[3] | proc_6_start_FIFO_blk[3] | proc_6_TLF_FIFO_blk[3] | proc_6_input_sync_blk[3] | proc_6_output_sync_blk[3]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_6_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_6_reg <= proc_dep_vld_vec_6;
        end
    end
    assign in_chan_dep_vld_vec_6[0] = dep_chan_vld_3_6;
    assign in_chan_dep_data_vec_6[16 : 0] = dep_chan_data_3_6;
    assign token_in_vec_6[0] = token_3_6;
    assign in_chan_dep_vld_vec_6[1] = dep_chan_vld_5_6;
    assign in_chan_dep_data_vec_6[33 : 17] = dep_chan_data_5_6;
    assign token_in_vec_6[1] = token_5_6;
    assign in_chan_dep_vld_vec_6[2] = dep_chan_vld_11_6;
    assign in_chan_dep_data_vec_6[50 : 34] = dep_chan_data_11_6;
    assign token_in_vec_6[2] = token_11_6;
    assign dep_chan_vld_6_5 = out_chan_dep_vld_vec_6[0];
    assign dep_chan_data_6_5 = out_chan_dep_data_6;
    assign token_6_5 = token_out_vec_6[0];
    assign dep_chan_vld_6_3 = out_chan_dep_vld_vec_6[1];
    assign dep_chan_data_6_3 = out_chan_dep_data_6;
    assign token_6_3 = token_out_vec_6[1];
    assign dep_chan_vld_6_11 = out_chan_dep_vld_vec_6[2];
    assign dep_chan_data_6_11 = out_chan_dep_data_6;
    assign token_6_11 = token_out_vec_6[2];
    assign dep_chan_vld_6_1 = out_chan_dep_vld_vec_6[3];
    assign dep_chan_data_6_1 = out_chan_dep_data_6;
    assign token_6_1 = token_out_vec_6[3];

    // Process: AESL_inst_top.ConvertWeightToStream_U0
    AESL_deadlock_detect_unit #(17, 7, 6, 6) AESL_deadlock_detect_unit_7 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_7),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_7),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_7),
        .token_in_vec(token_in_vec_7),
        .dl_detect_in(dl_detect_out),
        .origin(origin[7]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_7),
        .out_chan_dep_data(out_chan_dep_data_7),
        .token_out_vec(token_out_vec_7),
        .dl_detect_out(dl_in_vec[7]));

    assign proc_7_data_FIFO_blk[0] = 1'b0 | (~AESL_inst_top.ConvertWeightToStream_U0.grp_ConvertWeightToStream_Pipeline_VITIS_LOOP_229_1_VITIS_LOOP_232_2_VITIS_LOOP_234_s_fu_180.fifo_conv_w_0_blk_n) | (~AESL_inst_top.ConvertWeightToStream_U0.grp_ConvertWeightToStream_Pipeline_VITIS_LOOP_229_1_VITIS_LOOP_232_2_VITIS_LOOP_234_s_fu_180.fifo_conv_w_1_blk_n) | (~AESL_inst_top.ConvertWeightToStream_U0.grp_ConvertWeightToStream_Pipeline_VITIS_LOOP_229_1_VITIS_LOOP_232_2_VITIS_LOOP_234_s_fu_180.fifo_conv_w_2_blk_n) | (~AESL_inst_top.ConvertWeightToStream_U0.grp_ConvertWeightToStream_Pipeline_VITIS_LOOP_229_1_VITIS_LOOP_232_2_VITIS_LOOP_234_s_fu_180.fifo_conv_w_3_blk_n) | (~AESL_inst_top.ConvertWeightToStream_U0.mode_c69_blk_n);
    assign proc_7_data_PIPO_blk[0] = 1'b0;
    assign proc_7_start_FIFO_blk[0] = 1'b0;
    assign proc_7_TLF_FIFO_blk[0] = 1'b0;
    assign proc_7_input_sync_blk[0] = 1'b0;
    assign proc_7_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_7[0] = dl_detect_out ? proc_dep_vld_vec_7_reg[0] : (proc_7_data_FIFO_blk[0] | proc_7_data_PIPO_blk[0] | proc_7_start_FIFO_blk[0] | proc_7_TLF_FIFO_blk[0] | proc_7_input_sync_blk[0] | proc_7_output_sync_blk[0]);
    assign proc_7_data_FIFO_blk[1] = 1'b0 | (~AESL_inst_top.ConvertWeightToStream_U0.grp_ConvertWeightToStream_Pipeline_VITIS_LOOP_251_5_VITIS_LOOP_254_6_VITIS_LOOP_257_s_fu_168.fifo_mm_w_blk_n) | (~AESL_inst_top.ConvertWeightToStream_U0.mode_c68_blk_n);
    assign proc_7_data_PIPO_blk[1] = 1'b0;
    assign proc_7_start_FIFO_blk[1] = 1'b0;
    assign proc_7_TLF_FIFO_blk[1] = 1'b0;
    assign proc_7_input_sync_blk[1] = 1'b0;
    assign proc_7_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_7[1] = dl_detect_out ? proc_dep_vld_vec_7_reg[1] : (proc_7_data_FIFO_blk[1] | proc_7_data_PIPO_blk[1] | proc_7_start_FIFO_blk[1] | proc_7_TLF_FIFO_blk[1] | proc_7_input_sync_blk[1] | proc_7_output_sync_blk[1]);
    assign proc_7_data_FIFO_blk[2] = 1'b0;
    assign proc_7_data_PIPO_blk[2] = 1'b0;
    assign proc_7_start_FIFO_blk[2] = 1'b0;
    assign proc_7_TLF_FIFO_blk[2] = 1'b0;
    assign proc_7_input_sync_blk[2] = 1'b0 | (AESL_inst_top.ap_sync_ConvertWeightToStream_U0_ap_ready & AESL_inst_top.ConvertWeightToStream_U0.ap_idle & ~AESL_inst_top.ap_sync_entry_proc_U0_ap_ready);
    assign proc_7_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_7[2] = dl_detect_out ? proc_dep_vld_vec_7_reg[2] : (proc_7_data_FIFO_blk[2] | proc_7_data_PIPO_blk[2] | proc_7_start_FIFO_blk[2] | proc_7_TLF_FIFO_blk[2] | proc_7_input_sync_blk[2] | proc_7_output_sync_blk[2]);
    assign proc_7_data_FIFO_blk[3] = 1'b0;
    assign proc_7_data_PIPO_blk[3] = 1'b0;
    assign proc_7_start_FIFO_blk[3] = 1'b0;
    assign proc_7_TLF_FIFO_blk[3] = 1'b0;
    assign proc_7_input_sync_blk[3] = 1'b0 | (AESL_inst_top.ap_sync_ConvertWeightToStream_U0_ap_ready & AESL_inst_top.ConvertWeightToStream_U0.ap_idle & ~AESL_inst_top.ap_sync_Block_entry3_proc_U0_ap_ready);
    assign proc_7_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_7[3] = dl_detect_out ? proc_dep_vld_vec_7_reg[3] : (proc_7_data_FIFO_blk[3] | proc_7_data_PIPO_blk[3] | proc_7_start_FIFO_blk[3] | proc_7_TLF_FIFO_blk[3] | proc_7_input_sync_blk[3] | proc_7_output_sync_blk[3]);
    assign proc_7_data_FIFO_blk[4] = 1'b0;
    assign proc_7_data_PIPO_blk[4] = 1'b0;
    assign proc_7_start_FIFO_blk[4] = 1'b0;
    assign proc_7_TLF_FIFO_blk[4] = 1'b0;
    assign proc_7_input_sync_blk[4] = 1'b0 | (AESL_inst_top.ap_sync_ConvertWeightToStream_U0_ap_ready & AESL_inst_top.ConvertWeightToStream_U0.ap_idle & ~AESL_inst_top.ap_sync_ConvertBias_BN_U0_ap_ready);
    assign proc_7_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_7[4] = dl_detect_out ? proc_dep_vld_vec_7_reg[4] : (proc_7_data_FIFO_blk[4] | proc_7_data_PIPO_blk[4] | proc_7_start_FIFO_blk[4] | proc_7_TLF_FIFO_blk[4] | proc_7_input_sync_blk[4] | proc_7_output_sync_blk[4]);
    assign proc_7_data_FIFO_blk[5] = 1'b0;
    assign proc_7_data_PIPO_blk[5] = 1'b0;
    assign proc_7_start_FIFO_blk[5] = 1'b0;
    assign proc_7_TLF_FIFO_blk[5] = 1'b0;
    assign proc_7_input_sync_blk[5] = 1'b0 | (AESL_inst_top.ap_sync_ConvertWeightToStream_U0_ap_ready & AESL_inst_top.ConvertWeightToStream_U0.ap_idle & ~AESL_inst_top.ap_sync_ConvertInputToStream_U0_ap_ready);
    assign proc_7_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_7[5] = dl_detect_out ? proc_dep_vld_vec_7_reg[5] : (proc_7_data_FIFO_blk[5] | proc_7_data_PIPO_blk[5] | proc_7_start_FIFO_blk[5] | proc_7_TLF_FIFO_blk[5] | proc_7_input_sync_blk[5] | proc_7_output_sync_blk[5]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_7_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_7_reg <= proc_dep_vld_vec_7;
        end
    end
    assign in_chan_dep_vld_vec_7[0] = dep_chan_vld_0_7;
    assign in_chan_dep_data_vec_7[16 : 0] = dep_chan_data_0_7;
    assign token_in_vec_7[0] = token_0_7;
    assign in_chan_dep_vld_vec_7[1] = dep_chan_vld_1_7;
    assign in_chan_dep_data_vec_7[33 : 17] = dep_chan_data_1_7;
    assign token_in_vec_7[1] = token_1_7;
    assign in_chan_dep_vld_vec_7[2] = dep_chan_vld_2_7;
    assign in_chan_dep_data_vec_7[50 : 34] = dep_chan_data_2_7;
    assign token_in_vec_7[2] = token_2_7;
    assign in_chan_dep_vld_vec_7[3] = dep_chan_vld_3_7;
    assign in_chan_dep_data_vec_7[67 : 51] = dep_chan_data_3_7;
    assign token_in_vec_7[3] = token_3_7;
    assign in_chan_dep_vld_vec_7[4] = dep_chan_vld_8_7;
    assign in_chan_dep_data_vec_7[84 : 68] = dep_chan_data_8_7;
    assign token_in_vec_7[4] = token_8_7;
    assign in_chan_dep_vld_vec_7[5] = dep_chan_vld_9_7;
    assign in_chan_dep_data_vec_7[101 : 85] = dep_chan_data_9_7;
    assign token_in_vec_7[5] = token_9_7;
    assign dep_chan_vld_7_8 = out_chan_dep_vld_vec_7[0];
    assign dep_chan_data_7_8 = out_chan_dep_data_7;
    assign token_7_8 = token_out_vec_7[0];
    assign dep_chan_vld_7_9 = out_chan_dep_vld_vec_7[1];
    assign dep_chan_data_7_9 = out_chan_dep_data_7;
    assign token_7_9 = token_out_vec_7[1];
    assign dep_chan_vld_7_0 = out_chan_dep_vld_vec_7[2];
    assign dep_chan_data_7_0 = out_chan_dep_data_7;
    assign token_7_0 = token_out_vec_7[2];
    assign dep_chan_vld_7_1 = out_chan_dep_vld_vec_7[3];
    assign dep_chan_data_7_1 = out_chan_dep_data_7;
    assign token_7_1 = token_out_vec_7[3];
    assign dep_chan_vld_7_2 = out_chan_dep_vld_vec_7[4];
    assign dep_chan_data_7_2 = out_chan_dep_data_7;
    assign token_7_2 = token_out_vec_7[4];
    assign dep_chan_vld_7_3 = out_chan_dep_vld_vec_7[5];
    assign dep_chan_data_7_3 = out_chan_dep_data_7;
    assign token_7_3 = token_out_vec_7[5];

    // Process: AESL_inst_top.ConvWeightToArray_U0
    AESL_deadlock_detect_unit #(17, 8, 2, 3) AESL_deadlock_detect_unit_8 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_8),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_8),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_8),
        .token_in_vec(token_in_vec_8),
        .dl_detect_in(dl_detect_out),
        .origin(origin[8]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_8),
        .out_chan_dep_data(out_chan_dep_data_8),
        .token_out_vec(token_out_vec_8),
        .dl_detect_out(dl_in_vec[8]));

    assign proc_8_data_FIFO_blk[0] = 1'b0 | (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.fifo_conv_w_blk_n) | (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.fifo_conv_w_1_blk_n) | (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.fifo_conv_w_2_blk_n) | (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.fifo_conv_w_3_blk_n) | (~AESL_inst_top.ConvWeightToArray_U0.mode_blk_n);
    assign proc_8_data_PIPO_blk[0] = 1'b0;
    assign proc_8_start_FIFO_blk[0] = 1'b0;
    assign proc_8_TLF_FIFO_blk[0] = 1'b0;
    assign proc_8_input_sync_blk[0] = 1'b0;
    assign proc_8_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_8[0] = dl_detect_out ? proc_dep_vld_vec_8_reg[0] : (proc_8_data_FIFO_blk[0] | proc_8_data_PIPO_blk[0] | proc_8_start_FIFO_blk[0] | proc_8_TLF_FIFO_blk[0] | proc_8_input_sync_blk[0] | proc_8_output_sync_blk[0]);
    assign proc_8_data_FIFO_blk[1] = 1'b0 | (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.Conv_SA_W_blk_n) | (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.Conv_SA_W_1_blk_n) | (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.Conv_SA_W_2_blk_n) | (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.Conv_SA_W_3_blk_n) | (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.Conv_SA_W_4_blk_n) | (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.Conv_SA_W_5_blk_n) | (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.Conv_SA_W_6_blk_n) | (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.Conv_SA_W_7_blk_n) | (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.Conv_SA_W_8_blk_n) | (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.Conv_SA_W_9_blk_n) | (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.Conv_SA_W_10_blk_n) | (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.Conv_SA_W_11_blk_n) | (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.Conv_SA_W_12_blk_n) | (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.Conv_SA_W_13_blk_n) | (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.Conv_SA_W_14_blk_n) | (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.Conv_SA_W_15_blk_n) | (~AESL_inst_top.ConvWeightToArray_U0.num_w_sa_loc_c_blk_n) | (~AESL_inst_top.ConvWeightToArray_U0.mode_c67_blk_n);
    assign proc_8_data_PIPO_blk[1] = 1'b0;
    assign proc_8_start_FIFO_blk[1] = 1'b0 | (~AESL_inst_top.start_for_MuxWeightStream_U0_U.if_full_n & AESL_inst_top.ConvWeightToArray_U0.ap_start & ~AESL_inst_top.ConvWeightToArray_U0.real_start & (trans_in_cnt_1 == trans_out_cnt_1) & ~AESL_inst_top.start_for_MuxWeightStream_U0_U.if_read);
    assign proc_8_TLF_FIFO_blk[1] = 1'b0;
    assign proc_8_input_sync_blk[1] = 1'b0;
    assign proc_8_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_8[1] = dl_detect_out ? proc_dep_vld_vec_8_reg[1] : (proc_8_data_FIFO_blk[1] | proc_8_data_PIPO_blk[1] | proc_8_start_FIFO_blk[1] | proc_8_TLF_FIFO_blk[1] | proc_8_input_sync_blk[1] | proc_8_output_sync_blk[1]);
    assign proc_8_data_FIFO_blk[2] = 1'b0;
    assign proc_8_data_PIPO_blk[2] = 1'b0;
    assign proc_8_start_FIFO_blk[2] = 1'b0;
    assign proc_8_TLF_FIFO_blk[2] = 1'b0 | (~AESL_inst_top.num_w_sa_loc_c36_channel_U.if_empty_n & AESL_inst_top.ConvWeightToArray_U0.ap_idle & ~AESL_inst_top.num_w_sa_loc_c36_channel_U.if_write);
    assign proc_8_input_sync_blk[2] = 1'b0;
    assign proc_8_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_8[2] = dl_detect_out ? proc_dep_vld_vec_8_reg[2] : (proc_8_data_FIFO_blk[2] | proc_8_data_PIPO_blk[2] | proc_8_start_FIFO_blk[2] | proc_8_TLF_FIFO_blk[2] | proc_8_input_sync_blk[2] | proc_8_output_sync_blk[2]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_8_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_8_reg <= proc_dep_vld_vec_8;
        end
    end
    assign in_chan_dep_vld_vec_8[0] = dep_chan_vld_7_8;
    assign in_chan_dep_data_vec_8[16 : 0] = dep_chan_data_7_8;
    assign token_in_vec_8[0] = token_7_8;
    assign in_chan_dep_vld_vec_8[1] = dep_chan_vld_10_8;
    assign in_chan_dep_data_vec_8[33 : 17] = dep_chan_data_10_8;
    assign token_in_vec_8[1] = token_10_8;
    assign dep_chan_vld_8_7 = out_chan_dep_vld_vec_8[0];
    assign dep_chan_data_8_7 = out_chan_dep_data_8;
    assign token_8_7 = token_out_vec_8[0];
    assign dep_chan_vld_8_10 = out_chan_dep_vld_vec_8[1];
    assign dep_chan_data_8_10 = out_chan_dep_data_8;
    assign token_8_10 = token_out_vec_8[1];
    assign dep_chan_vld_8_1 = out_chan_dep_vld_vec_8[2];
    assign dep_chan_data_8_1 = out_chan_dep_data_8;
    assign token_8_1 = token_out_vec_8[2];

    // Process: AESL_inst_top.MMWeightToArray_U0
    AESL_deadlock_detect_unit #(17, 9, 2, 3) AESL_deadlock_detect_unit_9 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_9),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_9),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_9),
        .token_in_vec(token_in_vec_9),
        .dl_detect_in(dl_detect_out),
        .origin(origin[9]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_9),
        .out_chan_dep_data(out_chan_dep_data_9),
        .token_out_vec(token_out_vec_9),
        .dl_detect_out(dl_in_vec[9]));

    assign proc_9_data_FIFO_blk[0] = 1'b0 | (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.fifo_mm_w_blk_n) | (~AESL_inst_top.MMWeightToArray_U0.mode_blk_n);
    assign proc_9_data_PIPO_blk[0] = 1'b0;
    assign proc_9_start_FIFO_blk[0] = 1'b0;
    assign proc_9_TLF_FIFO_blk[0] = 1'b0;
    assign proc_9_input_sync_blk[0] = 1'b0;
    assign proc_9_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_9[0] = dl_detect_out ? proc_dep_vld_vec_9_reg[0] : (proc_9_data_FIFO_blk[0] | proc_9_data_PIPO_blk[0] | proc_9_start_FIFO_blk[0] | proc_9_TLF_FIFO_blk[0] | proc_9_input_sync_blk[0] | proc_9_output_sync_blk[0]);
    assign proc_9_data_FIFO_blk[1] = 1'b0 | (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.MM_SA_W_blk_n) | (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.MM_SA_W_1_blk_n) | (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.MM_SA_W_2_blk_n) | (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.MM_SA_W_3_blk_n) | (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.MM_SA_W_4_blk_n) | (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.MM_SA_W_5_blk_n) | (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.MM_SA_W_6_blk_n) | (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.MM_SA_W_7_blk_n) | (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.MM_SA_W_8_blk_n) | (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.MM_SA_W_9_blk_n) | (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.MM_SA_W_10_blk_n) | (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.MM_SA_W_11_blk_n) | (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.MM_SA_W_12_blk_n) | (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.MM_SA_W_13_blk_n) | (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.MM_SA_W_14_blk_n) | (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.MM_SA_W_15_blk_n);
    assign proc_9_data_PIPO_blk[1] = 1'b0;
    assign proc_9_start_FIFO_blk[1] = 1'b0;
    assign proc_9_TLF_FIFO_blk[1] = 1'b0;
    assign proc_9_input_sync_blk[1] = 1'b0;
    assign proc_9_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_9[1] = dl_detect_out ? proc_dep_vld_vec_9_reg[1] : (proc_9_data_FIFO_blk[1] | proc_9_data_PIPO_blk[1] | proc_9_start_FIFO_blk[1] | proc_9_TLF_FIFO_blk[1] | proc_9_input_sync_blk[1] | proc_9_output_sync_blk[1]);
    assign proc_9_data_FIFO_blk[2] = 1'b0;
    assign proc_9_data_PIPO_blk[2] = 1'b0;
    assign proc_9_start_FIFO_blk[2] = 1'b0;
    assign proc_9_TLF_FIFO_blk[2] = 1'b0 | (~AESL_inst_top.num_w_sa_loc_c35_channel_U.if_empty_n & AESL_inst_top.MMWeightToArray_U0.ap_idle & ~AESL_inst_top.num_w_sa_loc_c35_channel_U.if_write);
    assign proc_9_input_sync_blk[2] = 1'b0;
    assign proc_9_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_9[2] = dl_detect_out ? proc_dep_vld_vec_9_reg[2] : (proc_9_data_FIFO_blk[2] | proc_9_data_PIPO_blk[2] | proc_9_start_FIFO_blk[2] | proc_9_TLF_FIFO_blk[2] | proc_9_input_sync_blk[2] | proc_9_output_sync_blk[2]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_9_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_9_reg <= proc_dep_vld_vec_9;
        end
    end
    assign in_chan_dep_vld_vec_9[0] = dep_chan_vld_7_9;
    assign in_chan_dep_data_vec_9[16 : 0] = dep_chan_data_7_9;
    assign token_in_vec_9[0] = token_7_9;
    assign in_chan_dep_vld_vec_9[1] = dep_chan_vld_10_9;
    assign in_chan_dep_data_vec_9[33 : 17] = dep_chan_data_10_9;
    assign token_in_vec_9[1] = token_10_9;
    assign dep_chan_vld_9_7 = out_chan_dep_vld_vec_9[0];
    assign dep_chan_data_9_7 = out_chan_dep_data_9;
    assign token_9_7 = token_out_vec_9[0];
    assign dep_chan_vld_9_10 = out_chan_dep_vld_vec_9[1];
    assign dep_chan_data_9_10 = out_chan_dep_data_9;
    assign token_9_10 = token_out_vec_9[1];
    assign dep_chan_vld_9_1 = out_chan_dep_vld_vec_9[2];
    assign dep_chan_data_9_1 = out_chan_dep_data_9;
    assign token_9_1 = token_out_vec_9[2];

    // Process: AESL_inst_top.MuxWeightStream_U0
    AESL_deadlock_detect_unit #(17, 10, 3, 3) AESL_deadlock_detect_unit_10 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_10),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_10),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_10),
        .token_in_vec(token_in_vec_10),
        .dl_detect_in(dl_detect_out),
        .origin(origin[10]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_10),
        .out_chan_dep_data(out_chan_dep_data_10),
        .token_out_vec(token_out_vec_10),
        .dl_detect_out(dl_in_vec[10]));

    assign proc_10_data_FIFO_blk[0] = 1'b0 | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.Conv_SA_W_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.Conv_SA_W_1_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.Conv_SA_W_2_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.Conv_SA_W_3_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.Conv_SA_W_4_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.Conv_SA_W_5_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.Conv_SA_W_6_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.Conv_SA_W_7_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.Conv_SA_W_8_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.Conv_SA_W_9_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.Conv_SA_W_10_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.Conv_SA_W_11_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.Conv_SA_W_12_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.Conv_SA_W_13_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.Conv_SA_W_14_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.Conv_SA_W_15_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.num_w_sa_loc_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.mode_blk_n);
    assign proc_10_data_PIPO_blk[0] = 1'b0;
    assign proc_10_start_FIFO_blk[0] = 1'b0 | (~AESL_inst_top.start_for_MuxWeightStream_U0_U.if_empty_n & AESL_inst_top.MuxWeightStream_U0.ap_idle & ~AESL_inst_top.start_for_MuxWeightStream_U0_U.if_write);
    assign proc_10_TLF_FIFO_blk[0] = 1'b0;
    assign proc_10_input_sync_blk[0] = 1'b0;
    assign proc_10_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_10[0] = dl_detect_out ? proc_dep_vld_vec_10_reg[0] : (proc_10_data_FIFO_blk[0] | proc_10_data_PIPO_blk[0] | proc_10_start_FIFO_blk[0] | proc_10_TLF_FIFO_blk[0] | proc_10_input_sync_blk[0] | proc_10_output_sync_blk[0]);
    assign proc_10_data_FIFO_blk[1] = 1'b0 | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.MM_SA_W_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.MM_SA_W_1_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.MM_SA_W_2_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.MM_SA_W_3_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.MM_SA_W_4_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.MM_SA_W_5_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.MM_SA_W_6_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.MM_SA_W_7_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.MM_SA_W_8_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.MM_SA_W_9_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.MM_SA_W_10_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.MM_SA_W_11_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.MM_SA_W_12_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.MM_SA_W_13_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.MM_SA_W_14_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.MM_SA_W_15_blk_n);
    assign proc_10_data_PIPO_blk[1] = 1'b0;
    assign proc_10_start_FIFO_blk[1] = 1'b0;
    assign proc_10_TLF_FIFO_blk[1] = 1'b0;
    assign proc_10_input_sync_blk[1] = 1'b0;
    assign proc_10_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_10[1] = dl_detect_out ? proc_dep_vld_vec_10_reg[1] : (proc_10_data_FIFO_blk[1] | proc_10_data_PIPO_blk[1] | proc_10_start_FIFO_blk[1] | proc_10_TLF_FIFO_blk[1] | proc_10_input_sync_blk[1] | proc_10_output_sync_blk[1]);
    assign proc_10_data_FIFO_blk[2] = 1'b0 | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.fifo_SA_W_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.fifo_SA_W_1_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.fifo_SA_W_2_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.fifo_SA_W_3_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.fifo_SA_W_4_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.fifo_SA_W_5_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.fifo_SA_W_6_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.fifo_SA_W_7_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.fifo_SA_W_8_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.fifo_SA_W_9_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.fifo_SA_W_10_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.fifo_SA_W_11_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.fifo_SA_W_12_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.fifo_SA_W_13_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.fifo_SA_W_14_blk_n) | (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.fifo_SA_W_15_blk_n);
    assign proc_10_data_PIPO_blk[2] = 1'b0;
    assign proc_10_start_FIFO_blk[2] = 1'b0;
    assign proc_10_TLF_FIFO_blk[2] = 1'b0;
    assign proc_10_input_sync_blk[2] = 1'b0;
    assign proc_10_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_10[2] = dl_detect_out ? proc_dep_vld_vec_10_reg[2] : (proc_10_data_FIFO_blk[2] | proc_10_data_PIPO_blk[2] | proc_10_start_FIFO_blk[2] | proc_10_TLF_FIFO_blk[2] | proc_10_input_sync_blk[2] | proc_10_output_sync_blk[2]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_10_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_10_reg <= proc_dep_vld_vec_10;
        end
    end
    assign in_chan_dep_vld_vec_10[0] = dep_chan_vld_8_10;
    assign in_chan_dep_data_vec_10[16 : 0] = dep_chan_data_8_10;
    assign token_in_vec_10[0] = token_8_10;
    assign in_chan_dep_vld_vec_10[1] = dep_chan_vld_9_10;
    assign in_chan_dep_data_vec_10[33 : 17] = dep_chan_data_9_10;
    assign token_in_vec_10[1] = token_9_10;
    assign in_chan_dep_vld_vec_10[2] = dep_chan_vld_11_10;
    assign in_chan_dep_data_vec_10[50 : 34] = dep_chan_data_11_10;
    assign token_in_vec_10[2] = token_11_10;
    assign dep_chan_vld_10_8 = out_chan_dep_vld_vec_10[0];
    assign dep_chan_data_10_8 = out_chan_dep_data_10;
    assign token_10_8 = token_out_vec_10[0];
    assign dep_chan_vld_10_9 = out_chan_dep_vld_vec_10[1];
    assign dep_chan_data_10_9 = out_chan_dep_data_10;
    assign token_10_9 = token_out_vec_10[1];
    assign dep_chan_vld_10_11 = out_chan_dep_vld_vec_10[2];
    assign dep_chan_data_10_11 = out_chan_dep_data_10;
    assign token_10_11 = token_out_vec_10[2];

    // Process: AESL_inst_top.Compute_U0
    AESL_deadlock_detect_unit #(17, 11, 4, 5) AESL_deadlock_detect_unit_11 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_11),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_11),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_11),
        .token_in_vec(token_in_vec_11),
        .dl_detect_in(dl_detect_out),
        .origin(origin[11]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_11),
        .out_chan_dep_data(out_chan_dep_data_11),
        .token_out_vec(token_out_vec_11),
        .dl_detect_out(dl_in_vec[11]));

    assign proc_11_data_FIFO_blk[0] = 1'b0 | (~AESL_inst_top.Compute_U0.grp_PE_fu_278.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_A_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_300.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_A_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_322.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_A_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_344.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_A_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_366.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_A_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_388.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_A_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_410.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_A_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_432.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_A_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_454.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_A_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_476.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_A_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_498.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_A_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_520.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_A_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_542.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_A_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_564.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_A_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_586.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_A_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_608.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_A_0_0_blk_n) | (~AESL_inst_top.Compute_U0.num_a_sa_2_loc_blk_n) | (~AESL_inst_top.Compute_U0.mode_blk_n);
    assign proc_11_data_PIPO_blk[0] = 1'b0;
    assign proc_11_start_FIFO_blk[0] = 1'b0;
    assign proc_11_TLF_FIFO_blk[0] = 1'b0;
    assign proc_11_input_sync_blk[0] = 1'b0;
    assign proc_11_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_11[0] = dl_detect_out ? proc_dep_vld_vec_11_reg[0] : (proc_11_data_FIFO_blk[0] | proc_11_data_PIPO_blk[0] | proc_11_start_FIFO_blk[0] | proc_11_TLF_FIFO_blk[0] | proc_11_input_sync_blk[0] | proc_11_output_sync_blk[0]);
    assign proc_11_data_FIFO_blk[1] = 1'b0 | (~AESL_inst_top.Compute_U0.grp_PE_fu_278.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_W_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_300.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_W_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_322.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_W_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_344.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_W_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_366.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_W_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_388.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_W_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_410.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_W_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_432.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_W_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_454.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_W_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_476.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_W_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_498.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_W_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_520.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_W_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_542.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_W_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_564.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_W_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_586.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_W_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_608.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_W_0_0_blk_n);
    assign proc_11_data_PIPO_blk[1] = 1'b0;
    assign proc_11_start_FIFO_blk[1] = 1'b0;
    assign proc_11_TLF_FIFO_blk[1] = 1'b0;
    assign proc_11_input_sync_blk[1] = 1'b0;
    assign proc_11_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_11[1] = dl_detect_out ? proc_dep_vld_vec_11_reg[1] : (proc_11_data_FIFO_blk[1] | proc_11_data_PIPO_blk[1] | proc_11_start_FIFO_blk[1] | proc_11_TLF_FIFO_blk[1] | proc_11_input_sync_blk[1] | proc_11_output_sync_blk[1]);
    assign proc_11_data_FIFO_blk[2] = 1'b0 | (~AESL_inst_top.Compute_U0.grp_PE_fu_278.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_278.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_1_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_278.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_2_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_278.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_3_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_300.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_300.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_1_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_300.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_2_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_300.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_3_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_322.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_322.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_1_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_322.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_2_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_322.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_3_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_344.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_344.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_1_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_344.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_2_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_344.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_3_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_366.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_366.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_1_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_366.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_2_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_366.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_3_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_388.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_388.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_1_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_388.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_2_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_388.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_3_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_410.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_410.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_1_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_410.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_2_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_410.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_3_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_432.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_432.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_1_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_432.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_2_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_432.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_3_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_454.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_454.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_1_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_454.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_2_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_454.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_3_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_476.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_476.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_1_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_476.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_2_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_476.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_3_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_498.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_498.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_1_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_498.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_2_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_498.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_3_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_520.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_520.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_1_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_520.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_2_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_520.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_3_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_542.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_542.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_1_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_542.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_2_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_542.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_3_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_564.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_564.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_1_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_564.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_2_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_564.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_3_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_586.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_586.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_1_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_586.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_2_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_586.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_3_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_608.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_0_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_608.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_1_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_608.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_2_blk_n) | (~AESL_inst_top.Compute_U0.grp_PE_fu_608.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_3_blk_n) | (~AESL_inst_top.Compute_U0.num_a_sa_2_loc_c_blk_n) | (~AESL_inst_top.Compute_U0.mode_c65_blk_n);
    assign proc_11_data_PIPO_blk[2] = 1'b0;
    assign proc_11_start_FIFO_blk[2] = 1'b0;
    assign proc_11_TLF_FIFO_blk[2] = 1'b0;
    assign proc_11_input_sync_blk[2] = 1'b0;
    assign proc_11_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_11[2] = dl_detect_out ? proc_dep_vld_vec_11_reg[2] : (proc_11_data_FIFO_blk[2] | proc_11_data_PIPO_blk[2] | proc_11_start_FIFO_blk[2] | proc_11_TLF_FIFO_blk[2] | proc_11_input_sync_blk[2] | proc_11_output_sync_blk[2]);
    assign proc_11_data_FIFO_blk[3] = 1'b0;
    assign proc_11_data_PIPO_blk[3] = 1'b0;
    assign proc_11_start_FIFO_blk[3] = 1'b0;
    assign proc_11_TLF_FIFO_blk[3] = 1'b0 | (~AESL_inst_top.out_c_1_loc_c41_channel_U.if_empty_n & AESL_inst_top.Compute_U0.ap_idle & ~AESL_inst_top.out_c_1_loc_c41_channel_U.if_write);
    assign proc_11_input_sync_blk[3] = 1'b0;
    assign proc_11_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_11[3] = dl_detect_out ? proc_dep_vld_vec_11_reg[3] : (proc_11_data_FIFO_blk[3] | proc_11_data_PIPO_blk[3] | proc_11_start_FIFO_blk[3] | proc_11_TLF_FIFO_blk[3] | proc_11_input_sync_blk[3] | proc_11_output_sync_blk[3]);
    assign proc_11_data_FIFO_blk[4] = 1'b0 | (~AESL_inst_top.Compute_U0.out_c_1_loc_c40_blk_n);
    assign proc_11_data_PIPO_blk[4] = 1'b0;
    assign proc_11_start_FIFO_blk[4] = 1'b0;
    assign proc_11_TLF_FIFO_blk[4] = 1'b0;
    assign proc_11_input_sync_blk[4] = 1'b0;
    assign proc_11_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_11[4] = dl_detect_out ? proc_dep_vld_vec_11_reg[4] : (proc_11_data_FIFO_blk[4] | proc_11_data_PIPO_blk[4] | proc_11_start_FIFO_blk[4] | proc_11_TLF_FIFO_blk[4] | proc_11_input_sync_blk[4] | proc_11_output_sync_blk[4]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_11_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_11_reg <= proc_dep_vld_vec_11;
        end
    end
    assign in_chan_dep_vld_vec_11[0] = dep_chan_vld_6_11;
    assign in_chan_dep_data_vec_11[16 : 0] = dep_chan_data_6_11;
    assign token_in_vec_11[0] = token_6_11;
    assign in_chan_dep_vld_vec_11[1] = dep_chan_vld_10_11;
    assign in_chan_dep_data_vec_11[33 : 17] = dep_chan_data_10_11;
    assign token_in_vec_11[1] = token_10_11;
    assign in_chan_dep_vld_vec_11[2] = dep_chan_vld_12_11;
    assign in_chan_dep_data_vec_11[50 : 34] = dep_chan_data_12_11;
    assign token_in_vec_11[2] = token_12_11;
    assign in_chan_dep_vld_vec_11[3] = dep_chan_vld_13_11;
    assign in_chan_dep_data_vec_11[67 : 51] = dep_chan_data_13_11;
    assign token_in_vec_11[3] = token_13_11;
    assign dep_chan_vld_11_6 = out_chan_dep_vld_vec_11[0];
    assign dep_chan_data_11_6 = out_chan_dep_data_11;
    assign token_11_6 = token_out_vec_11[0];
    assign dep_chan_vld_11_10 = out_chan_dep_vld_vec_11[1];
    assign dep_chan_data_11_10 = out_chan_dep_data_11;
    assign token_11_10 = token_out_vec_11[1];
    assign dep_chan_vld_11_12 = out_chan_dep_vld_vec_11[2];
    assign dep_chan_data_11_12 = out_chan_dep_data_11;
    assign token_11_12 = token_out_vec_11[2];
    assign dep_chan_vld_11_1 = out_chan_dep_vld_vec_11[3];
    assign dep_chan_data_11_1 = out_chan_dep_data_11;
    assign token_11_1 = token_out_vec_11[3];
    assign dep_chan_vld_11_13 = out_chan_dep_vld_vec_11[4];
    assign dep_chan_data_11_13 = out_chan_dep_data_11;
    assign token_11_13 = token_out_vec_11[4];

    // Process: AESL_inst_top.ConvertToOutStream_U0
    AESL_deadlock_detect_unit #(17, 12, 4, 4) AESL_deadlock_detect_unit_12 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_12),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_12),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_12),
        .token_in_vec(token_in_vec_12),
        .dl_detect_in(dl_detect_out),
        .origin(origin[12]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_12),
        .out_chan_dep_data(out_chan_dep_data_12),
        .token_out_vec(token_out_vec_12),
        .dl_detect_out(dl_in_vec[12]));

    assign proc_12_data_FIFO_blk[0] = 1'b0 | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_1_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_2_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_3_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_4_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_5_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_6_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_7_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_8_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_9_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_10_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_11_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_12_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_13_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_14_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_15_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_16_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_17_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_18_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_19_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_20_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_21_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_22_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_23_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_24_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_25_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_26_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_27_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_28_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_29_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_30_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_31_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_32_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_33_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_34_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_35_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_36_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_37_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_38_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_39_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_40_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_41_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_42_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_43_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_44_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_45_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_46_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_47_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_48_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_49_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_50_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_51_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_52_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_53_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_54_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_55_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_56_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_57_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_58_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_59_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_60_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_61_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_62_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_63_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.num_a_sa_2_loc_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.mode_blk_n);
    assign proc_12_data_PIPO_blk[0] = 1'b0;
    assign proc_12_start_FIFO_blk[0] = 1'b0;
    assign proc_12_TLF_FIFO_blk[0] = 1'b0;
    assign proc_12_input_sync_blk[0] = 1'b0;
    assign proc_12_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_12[0] = dl_detect_out ? proc_dep_vld_vec_12_reg[0] : (proc_12_data_FIFO_blk[0] | proc_12_data_PIPO_blk[0] | proc_12_start_FIFO_blk[0] | proc_12_TLF_FIFO_blk[0] | proc_12_input_sync_blk[0] | proc_12_output_sync_blk[0]);
    assign proc_12_data_FIFO_blk[1] = 1'b0 | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_570_1_fu_464.fifo_CONV3_ACC_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_570_1_fu_464.fifo_CONV3_ACC_1_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_570_1_fu_464.fifo_CONV3_ACC_2_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_570_1_fu_464.fifo_CONV3_ACC_3_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_570_1_fu_464.fifo_CONV3_ACC_4_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_570_1_fu_464.fifo_CONV3_ACC_5_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_570_1_fu_464.fifo_CONV3_ACC_6_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_570_1_fu_464.fifo_CONV3_ACC_7_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_570_1_fu_464.fifo_CONV3_ACC_8_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_570_1_fu_464.fifo_CONV3_ACC_9_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_570_1_fu_464.fifo_CONV3_ACC_10_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_570_1_fu_464.fifo_CONV3_ACC_11_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_570_1_fu_464.fifo_CONV3_ACC_12_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_570_1_fu_464.fifo_CONV3_ACC_13_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_570_1_fu_464.fifo_CONV3_ACC_14_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_570_1_fu_464.fifo_CONV3_ACC_15_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.N_c_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.mode_c64_blk_n);
    assign proc_12_data_PIPO_blk[1] = 1'b0;
    assign proc_12_start_FIFO_blk[1] = 1'b0;
    assign proc_12_TLF_FIFO_blk[1] = 1'b0;
    assign proc_12_input_sync_blk[1] = 1'b0;
    assign proc_12_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_12[1] = dl_detect_out ? proc_dep_vld_vec_12_reg[1] : (proc_12_data_FIFO_blk[1] | proc_12_data_PIPO_blk[1] | proc_12_start_FIFO_blk[1] | proc_12_TLF_FIFO_blk[1] | proc_12_input_sync_blk[1] | proc_12_output_sync_blk[1]);
    assign proc_12_data_FIFO_blk[2] = 1'b0 | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.MM_OUT_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.MM_OUT_1_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.MM_OUT_2_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.MM_OUT_3_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.MM_OUT_4_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.MM_OUT_5_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.MM_OUT_6_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.MM_OUT_7_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.MM_OUT_8_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.MM_OUT_9_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.MM_OUT_10_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.MM_OUT_11_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.MM_OUT_12_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.MM_OUT_13_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.MM_OUT_14_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.MM_OUT_15_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.R_c_blk_n);
    assign proc_12_data_PIPO_blk[2] = 1'b0;
    assign proc_12_start_FIFO_blk[2] = 1'b0;
    assign proc_12_TLF_FIFO_blk[2] = 1'b0;
    assign proc_12_input_sync_blk[2] = 1'b0;
    assign proc_12_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_12[2] = dl_detect_out ? proc_dep_vld_vec_12_reg[2] : (proc_12_data_FIFO_blk[2] | proc_12_data_PIPO_blk[2] | proc_12_start_FIFO_blk[2] | proc_12_TLF_FIFO_blk[2] | proc_12_input_sync_blk[2] | proc_12_output_sync_blk[2]);
    assign proc_12_data_FIFO_blk[3] = 1'b0 | (~AESL_inst_top.ConvertToOutStream_U0.R_blk_n) | (~AESL_inst_top.ConvertToOutStream_U0.N_blk_n);
    assign proc_12_data_PIPO_blk[3] = 1'b0;
    assign proc_12_start_FIFO_blk[3] = 1'b0 | (~AESL_inst_top.start_for_ConvertToOutStream_U0_U.if_empty_n & AESL_inst_top.ConvertToOutStream_U0.ap_idle & ~AESL_inst_top.start_for_ConvertToOutStream_U0_U.if_write);
    assign proc_12_TLF_FIFO_blk[3] = 1'b0;
    assign proc_12_input_sync_blk[3] = 1'b0;
    assign proc_12_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_12[3] = dl_detect_out ? proc_dep_vld_vec_12_reg[3] : (proc_12_data_FIFO_blk[3] | proc_12_data_PIPO_blk[3] | proc_12_start_FIFO_blk[3] | proc_12_TLF_FIFO_blk[3] | proc_12_input_sync_blk[3] | proc_12_output_sync_blk[3]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_12_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_12_reg <= proc_dep_vld_vec_12;
        end
    end
    assign in_chan_dep_vld_vec_12[0] = dep_chan_vld_5_12;
    assign in_chan_dep_data_vec_12[16 : 0] = dep_chan_data_5_12;
    assign token_in_vec_12[0] = token_5_12;
    assign in_chan_dep_vld_vec_12[1] = dep_chan_vld_11_12;
    assign in_chan_dep_data_vec_12[33 : 17] = dep_chan_data_11_12;
    assign token_in_vec_12[1] = token_11_12;
    assign in_chan_dep_vld_vec_12[2] = dep_chan_vld_13_12;
    assign in_chan_dep_data_vec_12[50 : 34] = dep_chan_data_13_12;
    assign token_in_vec_12[2] = token_13_12;
    assign in_chan_dep_vld_vec_12[3] = dep_chan_vld_16_12;
    assign in_chan_dep_data_vec_12[67 : 51] = dep_chan_data_16_12;
    assign token_in_vec_12[3] = token_16_12;
    assign dep_chan_vld_12_11 = out_chan_dep_vld_vec_12[0];
    assign dep_chan_data_12_11 = out_chan_dep_data_12;
    assign token_12_11 = token_out_vec_12[0];
    assign dep_chan_vld_12_13 = out_chan_dep_vld_vec_12[1];
    assign dep_chan_data_12_13 = out_chan_dep_data_12;
    assign token_12_13 = token_out_vec_12[1];
    assign dep_chan_vld_12_16 = out_chan_dep_vld_vec_12[2];
    assign dep_chan_data_12_16 = out_chan_dep_data_12;
    assign token_12_16 = token_out_vec_12[2];
    assign dep_chan_vld_12_5 = out_chan_dep_vld_vec_12[3];
    assign dep_chan_data_12_5 = out_chan_dep_data_12;
    assign token_12_5 = token_out_vec_12[3];

    // Process: AESL_inst_top.ConvToOutStream_U0
    AESL_deadlock_detect_unit #(17, 13, 5, 6) AESL_deadlock_detect_unit_13 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_13),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_13),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_13),
        .token_in_vec(token_in_vec_13),
        .dl_detect_in(dl_detect_out),
        .origin(origin[13]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_13),
        .out_chan_dep_data(out_chan_dep_data_13),
        .token_out_vec(token_out_vec_13),
        .dl_detect_out(dl_in_vec[13]));

    assign proc_13_data_FIFO_blk[0] = 1'b0 | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.fifo_CONV3_ACC_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.fifo_CONV3_ACC_1_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.fifo_CONV3_ACC_2_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.fifo_CONV3_ACC_3_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.fifo_CONV3_ACC_4_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.fifo_CONV3_ACC_5_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.fifo_CONV3_ACC_6_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.fifo_CONV3_ACC_7_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.fifo_CONV3_ACC_8_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.fifo_CONV3_ACC_9_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.fifo_CONV3_ACC_10_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.fifo_CONV3_ACC_11_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.fifo_CONV3_ACC_12_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.fifo_CONV3_ACC_13_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.fifo_CONV3_ACC_14_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.fifo_CONV3_ACC_15_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.N_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.mode_blk_n);
    assign proc_13_data_PIPO_blk[0] = 1'b0;
    assign proc_13_start_FIFO_blk[0] = 1'b0;
    assign proc_13_TLF_FIFO_blk[0] = 1'b0;
    assign proc_13_input_sync_blk[0] = 1'b0;
    assign proc_13_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_13[0] = dl_detect_out ? proc_dep_vld_vec_13_reg[0] : (proc_13_data_FIFO_blk[0] | proc_13_data_PIPO_blk[0] | proc_13_start_FIFO_blk[0] | proc_13_TLF_FIFO_blk[0] | proc_13_input_sync_blk[0] | proc_13_output_sync_blk[0]);
    assign proc_13_data_FIFO_blk[1] = 1'b0 | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_1_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_2_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_3_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_4_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_5_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_6_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_7_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_8_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_9_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_10_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_11_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_12_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_13_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_14_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_15_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_16_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_17_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_18_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_19_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_20_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_21_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_22_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_23_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_24_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_25_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_26_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_27_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_28_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_29_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_30_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_31_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_32_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_33_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_34_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_35_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_36_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_37_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_38_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_39_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_40_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_41_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_42_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_43_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_44_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_45_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_46_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_47_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_48_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_49_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_50_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_51_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_52_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_53_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_54_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_55_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_56_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_57_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_58_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_59_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_60_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_61_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_62_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_63_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_64_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_65_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_66_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_67_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_68_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_69_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_70_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_71_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_72_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_73_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_74_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_75_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_76_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_77_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_78_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_79_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_80_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_81_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_82_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_83_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_84_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_85_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_86_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_87_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_88_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_89_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_90_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_91_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_92_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_93_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_94_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_95_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_96_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_97_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_98_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_99_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_100_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_101_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_102_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_103_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_104_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_105_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_106_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_107_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_108_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_109_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_110_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_111_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_112_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_113_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_114_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_115_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_116_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_117_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_118_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_119_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_120_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_121_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_122_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_123_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_124_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_125_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_126_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_127_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.out_r_1_loc_c37_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.out_c_1_loc_c39_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.M_c53_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.mode_c63_blk_n);
    assign proc_13_data_PIPO_blk[1] = 1'b0;
    assign proc_13_start_FIFO_blk[1] = 1'b0;
    assign proc_13_TLF_FIFO_blk[1] = 1'b0;
    assign proc_13_input_sync_blk[1] = 1'b0;
    assign proc_13_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_13[1] = dl_detect_out ? proc_dep_vld_vec_13_reg[1] : (proc_13_data_FIFO_blk[1] | proc_13_data_PIPO_blk[1] | proc_13_start_FIFO_blk[1] | proc_13_TLF_FIFO_blk[1] | proc_13_input_sync_blk[1] | proc_13_output_sync_blk[1]);
    assign proc_13_data_FIFO_blk[2] = 1'b0;
    assign proc_13_data_PIPO_blk[2] = 1'b0;
    assign proc_13_start_FIFO_blk[2] = 1'b0;
    assign proc_13_TLF_FIFO_blk[2] = 1'b0 | (~AESL_inst_top.out_r_1_loc_c38_channel_U.if_empty_n & AESL_inst_top.ConvToOutStream_U0.ap_idle & ~AESL_inst_top.out_r_1_loc_c38_channel_U.if_write);
    assign proc_13_input_sync_blk[2] = 1'b0;
    assign proc_13_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_13[2] = dl_detect_out ? proc_dep_vld_vec_13_reg[2] : (proc_13_data_FIFO_blk[2] | proc_13_data_PIPO_blk[2] | proc_13_start_FIFO_blk[2] | proc_13_TLF_FIFO_blk[2] | proc_13_input_sync_blk[2] | proc_13_output_sync_blk[2]);
    assign proc_13_data_FIFO_blk[3] = 1'b0 | (~AESL_inst_top.ConvToOutStream_U0.out_c_1_loc_blk_n);
    assign proc_13_data_PIPO_blk[3] = 1'b0;
    assign proc_13_start_FIFO_blk[3] = 1'b0;
    assign proc_13_TLF_FIFO_blk[3] = 1'b0;
    assign proc_13_input_sync_blk[3] = 1'b0;
    assign proc_13_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_13[3] = dl_detect_out ? proc_dep_vld_vec_13_reg[3] : (proc_13_data_FIFO_blk[3] | proc_13_data_PIPO_blk[3] | proc_13_start_FIFO_blk[3] | proc_13_TLF_FIFO_blk[3] | proc_13_input_sync_blk[3] | proc_13_output_sync_blk[3]);
    assign proc_13_data_FIFO_blk[4] = 1'b0 | (~AESL_inst_top.ConvToOutStream_U0.M_blk_n) | (~AESL_inst_top.ConvToOutStream_U0.K_blk_n);
    assign proc_13_data_PIPO_blk[4] = 1'b0;
    assign proc_13_start_FIFO_blk[4] = 1'b0;
    assign proc_13_TLF_FIFO_blk[4] = 1'b0;
    assign proc_13_input_sync_blk[4] = 1'b0;
    assign proc_13_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_13[4] = dl_detect_out ? proc_dep_vld_vec_13_reg[4] : (proc_13_data_FIFO_blk[4] | proc_13_data_PIPO_blk[4] | proc_13_start_FIFO_blk[4] | proc_13_TLF_FIFO_blk[4] | proc_13_input_sync_blk[4] | proc_13_output_sync_blk[4]);
    assign proc_13_data_FIFO_blk[5] = 1'b0 | (~AESL_inst_top.ConvToOutStream_U0.K_c_blk_n);
    assign proc_13_data_PIPO_blk[5] = 1'b0;
    assign proc_13_start_FIFO_blk[5] = 1'b0;
    assign proc_13_TLF_FIFO_blk[5] = 1'b0;
    assign proc_13_input_sync_blk[5] = 1'b0;
    assign proc_13_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_13[5] = dl_detect_out ? proc_dep_vld_vec_13_reg[5] : (proc_13_data_FIFO_blk[5] | proc_13_data_PIPO_blk[5] | proc_13_start_FIFO_blk[5] | proc_13_TLF_FIFO_blk[5] | proc_13_input_sync_blk[5] | proc_13_output_sync_blk[5]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_13_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_13_reg <= proc_dep_vld_vec_13;
        end
    end
    assign in_chan_dep_vld_vec_13[0] = dep_chan_vld_5_13;
    assign in_chan_dep_data_vec_13[16 : 0] = dep_chan_data_5_13;
    assign token_in_vec_13[0] = token_5_13;
    assign in_chan_dep_vld_vec_13[1] = dep_chan_vld_11_13;
    assign in_chan_dep_data_vec_13[33 : 17] = dep_chan_data_11_13;
    assign token_in_vec_13[1] = token_11_13;
    assign in_chan_dep_vld_vec_13[2] = dep_chan_vld_12_13;
    assign in_chan_dep_data_vec_13[50 : 34] = dep_chan_data_12_13;
    assign token_in_vec_13[2] = token_12_13;
    assign in_chan_dep_vld_vec_13[3] = dep_chan_vld_14_13;
    assign in_chan_dep_data_vec_13[67 : 51] = dep_chan_data_14_13;
    assign token_in_vec_13[3] = token_14_13;
    assign in_chan_dep_vld_vec_13[4] = dep_chan_vld_16_13;
    assign in_chan_dep_data_vec_13[84 : 68] = dep_chan_data_16_13;
    assign token_in_vec_13[4] = token_16_13;
    assign dep_chan_vld_13_12 = out_chan_dep_vld_vec_13[0];
    assign dep_chan_data_13_12 = out_chan_dep_data_13;
    assign token_13_12 = token_out_vec_13[0];
    assign dep_chan_vld_13_14 = out_chan_dep_vld_vec_13[1];
    assign dep_chan_data_13_14 = out_chan_dep_data_13;
    assign token_13_14 = token_out_vec_13[1];
    assign dep_chan_vld_13_1 = out_chan_dep_vld_vec_13[2];
    assign dep_chan_data_13_1 = out_chan_dep_data_13;
    assign token_13_1 = token_out_vec_13[2];
    assign dep_chan_vld_13_11 = out_chan_dep_vld_vec_13[3];
    assign dep_chan_data_13_11 = out_chan_dep_data_13;
    assign token_13_11 = token_out_vec_13[3];
    assign dep_chan_vld_13_5 = out_chan_dep_vld_vec_13[4];
    assign dep_chan_data_13_5 = out_chan_dep_data_13;
    assign token_13_5 = token_out_vec_13[4];
    assign dep_chan_vld_13_16 = out_chan_dep_vld_vec_13[5];
    assign dep_chan_data_13_16 = out_chan_dep_data_13;
    assign token_13_16 = token_out_vec_13[5];

    // Process: AESL_inst_top.ConvBias_U0
    AESL_deadlock_detect_unit #(17, 14, 3, 3) AESL_deadlock_detect_unit_14 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_14),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_14),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_14),
        .token_in_vec(token_in_vec_14),
        .dl_detect_in(dl_detect_out),
        .origin(origin[14]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_14),
        .out_chan_dep_data(out_chan_dep_data_14),
        .token_out_vec(token_out_vec_14),
        .dl_detect_out(dl_in_vec[14]));

    assign proc_14_data_FIFO_blk[0] = 1'b0 | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_1_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_2_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_3_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_4_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_5_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_6_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_7_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_8_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_9_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_10_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_11_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_12_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_13_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_14_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_15_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_16_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_17_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_18_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_19_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_20_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_21_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_22_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_23_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_24_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_25_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_26_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_27_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_28_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_29_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_30_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_31_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_32_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_33_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_34_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_35_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_36_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_37_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_38_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_39_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_40_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_41_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_42_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_43_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_44_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_45_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_46_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_47_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_48_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_49_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_50_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_51_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_52_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_53_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_54_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_55_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_56_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_57_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_58_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_59_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_60_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_61_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_62_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_63_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_64_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_65_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_66_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_67_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_68_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_69_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_70_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_71_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_72_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_73_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_74_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_75_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_76_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_77_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_78_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_79_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_80_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_81_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_82_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_83_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_84_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_85_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_86_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_87_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_88_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_89_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_90_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_91_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_92_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_93_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_94_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_95_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_96_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_97_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_98_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_99_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_100_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_101_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_102_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_103_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_104_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_105_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_106_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_107_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_108_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_109_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_110_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_111_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_112_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_113_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_114_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_115_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_116_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_117_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_118_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_119_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_120_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_121_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_122_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_123_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_124_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_125_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_126_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_127_blk_n) | (~AESL_inst_top.ConvBias_U0.out_r_1_loc_blk_n) | (~AESL_inst_top.ConvBias_U0.out_c_1_loc_blk_n) | (~AESL_inst_top.ConvBias_U0.M_blk_n) | (~AESL_inst_top.ConvBias_U0.mode_blk_n);
    assign proc_14_data_PIPO_blk[0] = 1'b0;
    assign proc_14_start_FIFO_blk[0] = 1'b0;
    assign proc_14_TLF_FIFO_blk[0] = 1'b0;
    assign proc_14_input_sync_blk[0] = 1'b0;
    assign proc_14_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_14[0] = dl_detect_out ? proc_dep_vld_vec_14_reg[0] : (proc_14_data_FIFO_blk[0] | proc_14_data_PIPO_blk[0] | proc_14_start_FIFO_blk[0] | proc_14_TLF_FIFO_blk[0] | proc_14_input_sync_blk[0] | proc_14_output_sync_blk[0]);
    assign proc_14_data_FIFO_blk[1] = 1'b0 | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_1_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_2_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_3_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_4_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_5_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_6_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_7_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_8_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_9_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_10_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_11_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_12_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_13_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_14_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_15_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_16_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_17_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_18_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_19_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_20_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_21_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_22_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_23_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_24_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_25_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_26_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_27_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_28_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_29_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_30_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_31_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_32_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_33_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_34_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_35_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_36_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_37_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_38_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_39_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_40_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_41_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_42_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_43_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_44_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_45_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_46_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_47_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_48_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_49_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_50_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_51_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_52_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_53_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_54_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_55_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_56_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_57_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_58_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_59_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_60_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_61_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_62_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_63_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_64_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_65_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_66_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_67_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_68_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_69_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_70_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_71_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_72_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_73_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_74_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_75_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_76_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_77_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_78_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_79_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_80_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_81_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_82_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_83_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_84_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_85_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_86_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_87_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_88_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_89_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_90_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_91_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_92_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_93_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_94_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_95_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_96_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_97_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_98_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_99_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_100_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_101_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_102_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_103_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_104_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_105_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_106_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_107_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_108_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_109_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_110_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_111_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_112_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_113_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_114_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_115_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_116_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_117_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_118_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_119_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_120_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_121_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_122_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_123_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_124_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_125_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_126_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_127_blk_n);
    assign proc_14_data_PIPO_blk[1] = 1'b0;
    assign proc_14_start_FIFO_blk[1] = 1'b0 | (~AESL_inst_top.start_for_ConvBias_U0_U.if_empty_n & AESL_inst_top.ConvBias_U0.ap_idle & ~AESL_inst_top.start_for_ConvBias_U0_U.if_write);
    assign proc_14_TLF_FIFO_blk[1] = 1'b0;
    assign proc_14_input_sync_blk[1] = 1'b0;
    assign proc_14_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_14[1] = dl_detect_out ? proc_dep_vld_vec_14_reg[1] : (proc_14_data_FIFO_blk[1] | proc_14_data_PIPO_blk[1] | proc_14_start_FIFO_blk[1] | proc_14_TLF_FIFO_blk[1] | proc_14_input_sync_blk[1] | proc_14_output_sync_blk[1]);
    assign proc_14_data_FIFO_blk[2] = 1'b0 | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_1_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_2_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_3_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_4_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_5_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_6_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_7_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_8_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_9_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_10_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_11_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_12_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_13_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_14_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_15_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_16_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_17_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_18_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_19_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_20_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_21_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_22_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_23_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_24_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_25_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_26_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_27_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_28_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_29_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_30_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_31_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_32_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_33_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_34_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_35_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_36_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_37_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_38_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_39_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_40_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_41_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_42_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_43_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_44_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_45_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_46_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_47_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_48_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_49_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_50_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_51_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_52_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_53_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_54_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_55_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_56_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_57_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_58_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_59_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_60_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_61_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_62_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_63_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_64_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_65_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_66_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_67_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_68_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_69_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_70_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_71_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_72_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_73_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_74_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_75_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_76_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_77_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_78_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_79_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_80_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_81_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_82_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_83_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_84_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_85_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_86_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_87_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_88_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_89_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_90_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_91_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_92_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_93_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_94_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_95_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_96_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_97_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_98_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_99_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_100_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_101_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_102_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_103_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_104_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_105_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_106_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_107_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_108_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_109_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_110_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_111_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_112_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_113_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_114_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_115_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_116_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_117_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_118_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_119_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_120_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_121_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_122_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_123_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_124_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_125_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_126_blk_n) | (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_127_blk_n) | (~AESL_inst_top.ConvBias_U0.out_r_1_loc_c_blk_n) | (~AESL_inst_top.ConvBias_U0.out_c_1_loc_c_blk_n) | (~AESL_inst_top.ConvBias_U0.M_c52_blk_n) | (~AESL_inst_top.ConvBias_U0.mode_c62_blk_n);
    assign proc_14_data_PIPO_blk[2] = 1'b0;
    assign proc_14_start_FIFO_blk[2] = 1'b0;
    assign proc_14_TLF_FIFO_blk[2] = 1'b0;
    assign proc_14_input_sync_blk[2] = 1'b0;
    assign proc_14_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_14[2] = dl_detect_out ? proc_dep_vld_vec_14_reg[2] : (proc_14_data_FIFO_blk[2] | proc_14_data_PIPO_blk[2] | proc_14_start_FIFO_blk[2] | proc_14_TLF_FIFO_blk[2] | proc_14_input_sync_blk[2] | proc_14_output_sync_blk[2]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_14_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_14_reg <= proc_dep_vld_vec_14;
        end
    end
    assign in_chan_dep_vld_vec_14[0] = dep_chan_vld_2_14;
    assign in_chan_dep_data_vec_14[16 : 0] = dep_chan_data_2_14;
    assign token_in_vec_14[0] = token_2_14;
    assign in_chan_dep_vld_vec_14[1] = dep_chan_vld_13_14;
    assign in_chan_dep_data_vec_14[33 : 17] = dep_chan_data_13_14;
    assign token_in_vec_14[1] = token_13_14;
    assign in_chan_dep_vld_vec_14[2] = dep_chan_vld_15_14;
    assign in_chan_dep_data_vec_14[50 : 34] = dep_chan_data_15_14;
    assign token_in_vec_14[2] = token_15_14;
    assign dep_chan_vld_14_13 = out_chan_dep_vld_vec_14[0];
    assign dep_chan_data_14_13 = out_chan_dep_data_14;
    assign token_14_13 = token_out_vec_14[0];
    assign dep_chan_vld_14_2 = out_chan_dep_vld_vec_14[1];
    assign dep_chan_data_14_2 = out_chan_dep_data_14;
    assign token_14_2 = token_out_vec_14[1];
    assign dep_chan_vld_14_15 = out_chan_dep_vld_vec_14[2];
    assign dep_chan_data_14_15 = out_chan_dep_data_14;
    assign token_14_15 = token_out_vec_14[2];

    // Process: AESL_inst_top.ConvBN_U0
    AESL_deadlock_detect_unit #(17, 15, 3, 3) AESL_deadlock_detect_unit_15 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_15),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_15),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_15),
        .token_in_vec(token_in_vec_15),
        .dl_detect_in(dl_detect_out),
        .origin(origin[15]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_15),
        .out_chan_dep_data(out_chan_dep_data_15),
        .token_out_vec(token_out_vec_15),
        .dl_detect_out(dl_in_vec[15]));

    assign proc_15_data_FIFO_blk[0] = 1'b0 | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_1_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_2_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_3_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_4_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_5_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_6_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_7_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_8_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_9_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_10_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_11_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_12_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_13_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_14_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_15_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_16_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_17_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_18_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_19_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_20_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_21_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_22_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_23_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_24_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_25_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_26_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_27_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_28_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_29_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_30_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_31_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_32_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_33_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_34_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_35_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_36_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_37_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_38_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_39_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_40_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_41_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_42_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_43_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_44_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_45_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_46_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_47_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_48_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_49_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_50_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_51_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_52_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_53_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_54_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_55_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_56_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_57_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_58_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_59_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_60_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_61_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_62_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_63_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_64_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_65_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_66_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_67_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_68_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_69_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_70_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_71_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_72_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_73_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_74_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_75_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_76_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_77_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_78_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_79_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_80_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_81_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_82_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_83_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_84_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_85_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_86_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_87_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_88_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_89_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_90_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_91_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_92_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_93_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_94_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_95_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_96_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_97_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_98_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_99_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_100_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_101_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_102_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_103_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_104_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_105_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_106_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_107_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_108_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_109_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_110_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_111_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_112_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_113_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_114_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_115_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_116_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_117_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_118_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_119_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_120_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_121_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_122_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_123_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_124_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_125_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_126_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_127_blk_n) | (~AESL_inst_top.ConvBN_U0.out_r_1_loc_blk_n) | (~AESL_inst_top.ConvBN_U0.out_c_1_loc_blk_n) | (~AESL_inst_top.ConvBN_U0.M_blk_n) | (~AESL_inst_top.ConvBN_U0.mode_blk_n);
    assign proc_15_data_PIPO_blk[0] = 1'b0;
    assign proc_15_start_FIFO_blk[0] = 1'b0;
    assign proc_15_TLF_FIFO_blk[0] = 1'b0;
    assign proc_15_input_sync_blk[0] = 1'b0;
    assign proc_15_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_15[0] = dl_detect_out ? proc_dep_vld_vec_15_reg[0] : (proc_15_data_FIFO_blk[0] | proc_15_data_PIPO_blk[0] | proc_15_start_FIFO_blk[0] | proc_15_TLF_FIFO_blk[0] | proc_15_input_sync_blk[0] | proc_15_output_sync_blk[0]);
    assign proc_15_data_FIFO_blk[1] = 1'b0 | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_1_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_2_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_3_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_4_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_5_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_6_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_7_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_8_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_9_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_10_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_11_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_12_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_13_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_14_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_15_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_16_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_17_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_18_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_19_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_20_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_21_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_22_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_23_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_24_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_25_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_26_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_27_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_28_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_29_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_30_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_31_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_32_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_33_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_34_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_35_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_36_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_37_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_38_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_39_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_40_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_41_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_42_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_43_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_44_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_45_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_46_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_47_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_48_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_49_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_50_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_51_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_52_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_53_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_54_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_55_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_56_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_57_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_58_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_59_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_60_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_61_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_62_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_63_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_64_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_65_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_66_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_67_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_68_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_69_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_70_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_71_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_72_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_73_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_74_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_75_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_76_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_77_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_78_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_79_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_80_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_81_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_82_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_83_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_84_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_85_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_86_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_87_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_88_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_89_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_90_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_91_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_92_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_93_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_94_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_95_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_96_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_97_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_98_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_99_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_100_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_101_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_102_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_103_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_104_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_105_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_106_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_107_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_108_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_109_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_110_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_111_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_112_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_113_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_114_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_115_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_116_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_117_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_118_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_119_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_120_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_121_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_122_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_123_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_124_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_125_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_126_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_127_blk_n) | (~AESL_inst_top.ConvBN_U0.M_c_blk_n) | (~AESL_inst_top.ConvBN_U0.mode_c_blk_n);
    assign proc_15_data_PIPO_blk[1] = 1'b0;
    assign proc_15_start_FIFO_blk[1] = 1'b0;
    assign proc_15_TLF_FIFO_blk[1] = 1'b0;
    assign proc_15_input_sync_blk[1] = 1'b0;
    assign proc_15_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_15[1] = dl_detect_out ? proc_dep_vld_vec_15_reg[1] : (proc_15_data_FIFO_blk[1] | proc_15_data_PIPO_blk[1] | proc_15_start_FIFO_blk[1] | proc_15_TLF_FIFO_blk[1] | proc_15_input_sync_blk[1] | proc_15_output_sync_blk[1]);
    assign proc_15_data_FIFO_blk[2] = 1'b0 | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_1_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_2_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_3_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_4_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_5_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_6_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_7_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_8_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_9_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_10_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_11_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_12_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_13_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_14_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_15_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_16_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_17_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_18_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_19_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_20_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_21_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_22_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_23_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_24_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_25_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_26_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_27_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_28_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_29_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_30_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_31_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_32_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_33_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_34_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_35_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_36_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_37_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_38_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_39_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_40_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_41_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_42_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_43_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_44_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_45_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_46_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_47_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_48_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_49_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_50_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_51_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_52_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_53_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_54_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_55_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_56_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_57_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_58_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_59_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_60_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_61_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_62_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_63_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_64_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_65_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_66_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_67_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_68_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_69_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_70_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_71_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_72_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_73_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_74_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_75_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_76_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_77_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_78_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_79_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_80_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_81_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_82_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_83_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_84_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_85_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_86_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_87_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_88_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_89_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_90_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_91_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_92_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_93_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_94_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_95_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_96_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_97_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_98_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_99_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_100_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_101_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_102_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_103_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_104_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_105_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_106_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_107_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_108_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_109_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_110_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_111_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_112_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_113_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_114_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_115_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_116_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_117_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_118_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_119_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_120_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_121_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_122_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_123_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_124_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_125_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_126_blk_n) | (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_127_blk_n);
    assign proc_15_data_PIPO_blk[2] = 1'b0;
    assign proc_15_start_FIFO_blk[2] = 1'b0 | (~AESL_inst_top.start_for_ConvBN_U0_U.if_empty_n & AESL_inst_top.ConvBN_U0.ap_idle & ~AESL_inst_top.start_for_ConvBN_U0_U.if_write);
    assign proc_15_TLF_FIFO_blk[2] = 1'b0;
    assign proc_15_input_sync_blk[2] = 1'b0;
    assign proc_15_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_15[2] = dl_detect_out ? proc_dep_vld_vec_15_reg[2] : (proc_15_data_FIFO_blk[2] | proc_15_data_PIPO_blk[2] | proc_15_start_FIFO_blk[2] | proc_15_TLF_FIFO_blk[2] | proc_15_input_sync_blk[2] | proc_15_output_sync_blk[2]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_15_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_15_reg <= proc_dep_vld_vec_15;
        end
    end
    assign in_chan_dep_vld_vec_15[0] = dep_chan_vld_2_15;
    assign in_chan_dep_data_vec_15[16 : 0] = dep_chan_data_2_15;
    assign token_in_vec_15[0] = token_2_15;
    assign in_chan_dep_vld_vec_15[1] = dep_chan_vld_14_15;
    assign in_chan_dep_data_vec_15[33 : 17] = dep_chan_data_14_15;
    assign token_in_vec_15[1] = token_14_15;
    assign in_chan_dep_vld_vec_15[2] = dep_chan_vld_16_15;
    assign in_chan_dep_data_vec_15[50 : 34] = dep_chan_data_16_15;
    assign token_in_vec_15[2] = token_16_15;
    assign dep_chan_vld_15_14 = out_chan_dep_vld_vec_15[0];
    assign dep_chan_data_15_14 = out_chan_dep_data_15;
    assign token_15_14 = token_out_vec_15[0];
    assign dep_chan_vld_15_16 = out_chan_dep_vld_vec_15[1];
    assign dep_chan_data_15_16 = out_chan_dep_data_15;
    assign token_15_16 = token_out_vec_15[1];
    assign dep_chan_vld_15_2 = out_chan_dep_vld_vec_15[2];
    assign dep_chan_data_15_2 = out_chan_dep_data_15;
    assign token_15_2 = token_out_vec_15[2];

    // Process: AESL_inst_top.ResOutput_U0
    AESL_deadlock_detect_unit #(17, 16, 5, 5) AESL_deadlock_detect_unit_16 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_16),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_16),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_16),
        .token_in_vec(token_in_vec_16),
        .dl_detect_in(dl_detect_out),
        .origin(origin[16]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_16),
        .out_chan_dep_data(out_chan_dep_data_16),
        .token_out_vec(token_out_vec_16),
        .dl_detect_out(dl_in_vec[16]));

    assign proc_16_data_FIFO_blk[0] = 1'b0 | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_0_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_1_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_2_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_3_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_4_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_5_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_6_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_7_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_8_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_9_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_10_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_11_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_12_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_13_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_14_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_15_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_16_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_17_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_18_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_19_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_20_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_21_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_22_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_23_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_24_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_25_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_26_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_27_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_28_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_29_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_30_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_31_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_32_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_33_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_34_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_35_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_36_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_37_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_38_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_39_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_40_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_41_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_42_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_43_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_44_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_45_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_46_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_47_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_48_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_49_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_50_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_51_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_52_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_53_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_54_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_55_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_56_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_57_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_58_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_59_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_60_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_61_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_62_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_63_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_64_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_65_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_66_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_67_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_68_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_69_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_70_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_71_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_72_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_73_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_74_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_75_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_76_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_77_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_78_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_79_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_80_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_81_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_82_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_83_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_84_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_85_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_86_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_87_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_88_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_89_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_90_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_91_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_92_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_93_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_94_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_95_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_96_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_97_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_98_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_99_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_100_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_101_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_102_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_103_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_104_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_105_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_106_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_107_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_108_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_109_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_110_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_111_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_112_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_113_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_114_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_115_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_116_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_117_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_118_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_119_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_120_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_121_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_122_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_123_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_124_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_125_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_126_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_127_blk_n) | (~AESL_inst_top.ResOutput_U0.M_blk_n) | (~AESL_inst_top.ResOutput_U0.mode_blk_n);
    assign proc_16_data_PIPO_blk[0] = 1'b0;
    assign proc_16_start_FIFO_blk[0] = 1'b0;
    assign proc_16_TLF_FIFO_blk[0] = 1'b0;
    assign proc_16_input_sync_blk[0] = 1'b0;
    assign proc_16_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_16[0] = dl_detect_out ? proc_dep_vld_vec_16_reg[0] : (proc_16_data_FIFO_blk[0] | proc_16_data_PIPO_blk[0] | proc_16_start_FIFO_blk[0] | proc_16_TLF_FIFO_blk[0] | proc_16_input_sync_blk[0] | proc_16_output_sync_blk[0]);
    assign proc_16_data_FIFO_blk[1] = 1'b0 | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_734_4_VITIS_LOOP_737_5_VITIS_LOOP_740_6_VITIS_LOOP_fu_406.MM_OUT_0_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_734_4_VITIS_LOOP_737_5_VITIS_LOOP_740_6_VITIS_LOOP_fu_406.MM_OUT_1_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_734_4_VITIS_LOOP_737_5_VITIS_LOOP_740_6_VITIS_LOOP_fu_406.MM_OUT_2_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_734_4_VITIS_LOOP_737_5_VITIS_LOOP_740_6_VITIS_LOOP_fu_406.MM_OUT_3_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_734_4_VITIS_LOOP_737_5_VITIS_LOOP_740_6_VITIS_LOOP_fu_406.MM_OUT_4_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_734_4_VITIS_LOOP_737_5_VITIS_LOOP_740_6_VITIS_LOOP_fu_406.MM_OUT_5_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_734_4_VITIS_LOOP_737_5_VITIS_LOOP_740_6_VITIS_LOOP_fu_406.MM_OUT_6_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_734_4_VITIS_LOOP_737_5_VITIS_LOOP_740_6_VITIS_LOOP_fu_406.MM_OUT_7_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_734_4_VITIS_LOOP_737_5_VITIS_LOOP_740_6_VITIS_LOOP_fu_406.MM_OUT_8_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_734_4_VITIS_LOOP_737_5_VITIS_LOOP_740_6_VITIS_LOOP_fu_406.MM_OUT_9_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_734_4_VITIS_LOOP_737_5_VITIS_LOOP_740_6_VITIS_LOOP_fu_406.MM_OUT_10_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_734_4_VITIS_LOOP_737_5_VITIS_LOOP_740_6_VITIS_LOOP_fu_406.MM_OUT_11_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_734_4_VITIS_LOOP_737_5_VITIS_LOOP_740_6_VITIS_LOOP_fu_406.MM_OUT_12_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_734_4_VITIS_LOOP_737_5_VITIS_LOOP_740_6_VITIS_LOOP_fu_406.MM_OUT_13_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_734_4_VITIS_LOOP_737_5_VITIS_LOOP_740_6_VITIS_LOOP_fu_406.MM_OUT_14_blk_n) | (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_734_4_VITIS_LOOP_737_5_VITIS_LOOP_740_6_VITIS_LOOP_fu_406.MM_OUT_15_blk_n) | (~AESL_inst_top.ResOutput_U0.R_blk_n);
    assign proc_16_data_PIPO_blk[1] = 1'b0;
    assign proc_16_start_FIFO_blk[1] = 1'b0;
    assign proc_16_TLF_FIFO_blk[1] = 1'b0;
    assign proc_16_input_sync_blk[1] = 1'b0;
    assign proc_16_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_16[1] = dl_detect_out ? proc_dep_vld_vec_16_reg[1] : (proc_16_data_FIFO_blk[1] | proc_16_data_PIPO_blk[1] | proc_16_start_FIFO_blk[1] | proc_16_TLF_FIFO_blk[1] | proc_16_input_sync_blk[1] | proc_16_output_sync_blk[1]);
    assign proc_16_data_FIFO_blk[2] = 1'b0 | (~AESL_inst_top.ResOutput_U0.output_r_blk_n);
    assign proc_16_data_PIPO_blk[2] = 1'b0;
    assign proc_16_start_FIFO_blk[2] = 1'b0 | (~AESL_inst_top.start_for_ResOutput_U0_U.if_empty_n & AESL_inst_top.ResOutput_U0.ap_idle & ~AESL_inst_top.start_for_ResOutput_U0_U.if_write);
    assign proc_16_TLF_FIFO_blk[2] = 1'b0;
    assign proc_16_input_sync_blk[2] = 1'b0;
    assign proc_16_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_16[2] = dl_detect_out ? proc_dep_vld_vec_16_reg[2] : (proc_16_data_FIFO_blk[2] | proc_16_data_PIPO_blk[2] | proc_16_start_FIFO_blk[2] | proc_16_TLF_FIFO_blk[2] | proc_16_input_sync_blk[2] | proc_16_output_sync_blk[2]);
    assign proc_16_data_FIFO_blk[3] = 1'b0 | (~AESL_inst_top.ResOutput_U0.C_blk_n) | (~AESL_inst_top.ResOutput_U0.P_blk_n) | (~AESL_inst_top.ResOutput_U0.S_blk_n);
    assign proc_16_data_PIPO_blk[3] = 1'b0;
    assign proc_16_start_FIFO_blk[3] = 1'b0;
    assign proc_16_TLF_FIFO_blk[3] = 1'b0;
    assign proc_16_input_sync_blk[3] = 1'b0;
    assign proc_16_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_16[3] = dl_detect_out ? proc_dep_vld_vec_16_reg[3] : (proc_16_data_FIFO_blk[3] | proc_16_data_PIPO_blk[3] | proc_16_start_FIFO_blk[3] | proc_16_TLF_FIFO_blk[3] | proc_16_input_sync_blk[3] | proc_16_output_sync_blk[3]);
    assign proc_16_data_FIFO_blk[4] = 1'b0 | (~AESL_inst_top.ResOutput_U0.K_blk_n);
    assign proc_16_data_PIPO_blk[4] = 1'b0;
    assign proc_16_start_FIFO_blk[4] = 1'b0;
    assign proc_16_TLF_FIFO_blk[4] = 1'b0;
    assign proc_16_input_sync_blk[4] = 1'b0;
    assign proc_16_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_16[4] = dl_detect_out ? proc_dep_vld_vec_16_reg[4] : (proc_16_data_FIFO_blk[4] | proc_16_data_PIPO_blk[4] | proc_16_start_FIFO_blk[4] | proc_16_TLF_FIFO_blk[4] | proc_16_input_sync_blk[4] | proc_16_output_sync_blk[4]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_16_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_16_reg <= proc_dep_vld_vec_16;
        end
    end
    assign in_chan_dep_vld_vec_16[0] = dep_chan_vld_0_16;
    assign in_chan_dep_data_vec_16[16 : 0] = dep_chan_data_0_16;
    assign token_in_vec_16[0] = token_0_16;
    assign in_chan_dep_vld_vec_16[1] = dep_chan_vld_5_16;
    assign in_chan_dep_data_vec_16[33 : 17] = dep_chan_data_5_16;
    assign token_in_vec_16[1] = token_5_16;
    assign in_chan_dep_vld_vec_16[2] = dep_chan_vld_12_16;
    assign in_chan_dep_data_vec_16[50 : 34] = dep_chan_data_12_16;
    assign token_in_vec_16[2] = token_12_16;
    assign in_chan_dep_vld_vec_16[3] = dep_chan_vld_13_16;
    assign in_chan_dep_data_vec_16[67 : 51] = dep_chan_data_13_16;
    assign token_in_vec_16[3] = token_13_16;
    assign in_chan_dep_vld_vec_16[4] = dep_chan_vld_15_16;
    assign in_chan_dep_data_vec_16[84 : 68] = dep_chan_data_15_16;
    assign token_in_vec_16[4] = token_15_16;
    assign dep_chan_vld_16_15 = out_chan_dep_vld_vec_16[0];
    assign dep_chan_data_16_15 = out_chan_dep_data_16;
    assign token_16_15 = token_out_vec_16[0];
    assign dep_chan_vld_16_12 = out_chan_dep_vld_vec_16[1];
    assign dep_chan_data_16_12 = out_chan_dep_data_16;
    assign token_16_12 = token_out_vec_16[1];
    assign dep_chan_vld_16_0 = out_chan_dep_vld_vec_16[2];
    assign dep_chan_data_16_0 = out_chan_dep_data_16;
    assign token_16_0 = token_out_vec_16[2];
    assign dep_chan_vld_16_5 = out_chan_dep_vld_vec_16[3];
    assign dep_chan_data_16_5 = out_chan_dep_data_16;
    assign token_16_5 = token_out_vec_16[3];
    assign dep_chan_vld_16_13 = out_chan_dep_vld_vec_16[4];
    assign dep_chan_data_16_13 = out_chan_dep_data_16;
    assign token_16_13 = token_out_vec_16[4];


    wire [16:0] dl_in_vec_comb = dl_in_vec & ~{16{all_finish}};
    AESL_deadlock_report_unit #(17) AESL_deadlock_report_unit_inst (
        .dl_reset(dl_reset),
        .dl_clock(dl_clock),
        .dl_in_vec(dl_in_vec_comb),
        .trans_in_cnt_0(trans_in_cnt_0),
        .trans_out_cnt_0(trans_out_cnt_0),
        .trans_in_cnt_1(trans_in_cnt_1),
        .trans_out_cnt_1(trans_out_cnt_1),
        .trans_in_cnt_2(trans_in_cnt_2),
        .trans_out_cnt_2(trans_out_cnt_2),
        .trans_in_cnt_3(trans_in_cnt_3),
        .trans_out_cnt_3(trans_out_cnt_3),
        .ap_done_reg_0(ap_done_reg_0),
        .ap_done_reg_1(ap_done_reg_1),
        .ap_done_reg_2(ap_done_reg_2),
        .ap_done_reg_3(ap_done_reg_3),
        .ap_done_reg_4(ap_done_reg_4),
        .dl_detect_out(dl_detect_out),
        .origin(origin),
        .token_clear(token_clear));

endmodule
