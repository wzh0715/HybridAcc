`timescale 1 ns / 1 ps

module AESL_deadlock_report_unit #( parameter PROC_NUM = 4 ) (
    input dl_reset,
    input dl_clock,
    input [PROC_NUM - 1:0] dl_in_vec,
    input [15:0] trans_in_cnt_0,
    input [15:0] trans_out_cnt_0,
    input [15:0] trans_in_cnt_1,
    input [15:0] trans_out_cnt_1,
    input [15:0] trans_in_cnt_2,
    input [15:0] trans_out_cnt_2,
    input [15:0] trans_in_cnt_3,
    input [15:0] trans_out_cnt_3,
    input ap_done_reg_0,
    input ap_done_reg_1,
    input ap_done_reg_2,
    input ap_done_reg_3,
    input ap_done_reg_4,
    output dl_detect_out,
    output reg [PROC_NUM - 1:0] origin,
    output token_clear);
   
    // FSM states
    localparam ST_IDLE = 3'b000;
    localparam ST_FILTER_FAKE = 3'b001;
    localparam ST_DL_DETECTED = 3'b010;
    localparam ST_DL_REPORT = 3'b100;

    reg find_df_deadlock;
    reg [2:0] CS_fsm;
    reg [2:0] NS_fsm;
    reg [PROC_NUM - 1:0] dl_detect_reg;
    reg [PROC_NUM - 1:0] dl_done_reg;
    reg [PROC_NUM - 1:0] origin_reg;
    reg [PROC_NUM - 1:0] dl_in_vec_reg;
    reg [31:0] dl_keep_cnt;
    integer i;
    integer fp;

    // FSM State machine
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            CS_fsm <= ST_IDLE;
        end
        else begin
            CS_fsm <= NS_fsm;
        end
    end
    always @ (CS_fsm or dl_in_vec or dl_detect_reg or dl_done_reg or dl_in_vec or origin_reg or dl_keep_cnt) begin
        case (CS_fsm)
            ST_IDLE : begin
                if (|dl_in_vec) begin
                    NS_fsm = ST_FILTER_FAKE;
                end
                else begin
                    NS_fsm = ST_IDLE;
                end
            end
            ST_FILTER_FAKE: begin
                if (dl_keep_cnt >= 32'd1000) begin
                    NS_fsm = ST_DL_DETECTED;
                end
                else if (dl_detect_reg != (dl_detect_reg & dl_in_vec)) begin
                    NS_fsm = ST_IDLE;
                end
                else begin
                    NS_fsm = ST_FILTER_FAKE;
                end
            end
            ST_DL_DETECTED: begin
                // has unreported deadlock cycle
                if (dl_detect_reg != dl_done_reg) begin
                    NS_fsm = ST_DL_REPORT;
                end
                else begin
                    NS_fsm = ST_DL_DETECTED;
                end
            end
            ST_DL_REPORT: begin
                if (|(dl_in_vec & origin_reg)) begin
                    NS_fsm = ST_DL_DETECTED;
                end
                else begin
                    NS_fsm = ST_DL_REPORT;
                end
            end
            default: NS_fsm = ST_IDLE;
        endcase
    end

    // dl_detect_reg record the procs that first detect deadlock
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_detect_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_IDLE) begin
                dl_detect_reg <= dl_in_vec;
            end
        end
    end

    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_keep_cnt <= 32'h0;
        end
        else begin
            if (CS_fsm == ST_FILTER_FAKE && (dl_detect_reg == (dl_detect_reg & dl_in_vec))) begin
                dl_keep_cnt <= dl_keep_cnt + 32'h1;
            end
            else if (CS_fsm == ST_FILTER_FAKE && (dl_detect_reg != (dl_detect_reg & dl_in_vec))) begin
                dl_keep_cnt <= 32'h0;
            end
        end
    end

    // dl_detect_out keeps in high after deadlock detected
    assign dl_detect_out = (|dl_detect_reg) && (CS_fsm == ST_DL_DETECTED || CS_fsm == ST_DL_REPORT);

    // dl_done_reg record the cycles has been reported
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_done_reg <= 'b0;
        end
        else begin
            if ((CS_fsm == ST_DL_REPORT) && (|(dl_in_vec & dl_detect_reg) == 'b1)) begin
                dl_done_reg <= dl_done_reg | dl_in_vec;
            end
        end
    end

    // clear token once a cycle is done
    assign token_clear = (CS_fsm == ST_DL_REPORT) ? ((|(dl_in_vec & origin_reg)) ? 'b1 : 'b0) : 'b0;

    // origin_reg record the current cycle start id
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            origin_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED) begin
                origin_reg <= origin;
            end
        end
    end
   
    // origin will be valid for only one cycle
    wire [PROC_NUM*PROC_NUM - 1:0] origin_tmp;
    assign origin_tmp[PROC_NUM - 1:0] = (dl_detect_reg[0] & ~dl_done_reg[0]) ? 'b1 : 'b0;
    genvar j;
    generate
    for(j = 1;j < PROC_NUM;j = j + 1) begin: F1
        assign origin_tmp[j*PROC_NUM +: PROC_NUM] = (dl_detect_reg[j] & ~dl_done_reg[j]) ? ('b1 << j) : origin_tmp[(j - 1)*PROC_NUM +: PROC_NUM];
    end
    endgenerate
    always @ (CS_fsm or origin_tmp) begin
        if (CS_fsm == ST_DL_DETECTED) begin
            origin = origin_tmp[(PROC_NUM - 1)*PROC_NUM +: PROC_NUM];
        end
        else begin
            origin = 'b0;
        end
    end

    
    // dl_in_vec_reg record the current cycle dl_in_vec
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_in_vec_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED) begin
                dl_in_vec_reg <= origin;
            end
            else if (CS_fsm == ST_DL_REPORT) begin
                dl_in_vec_reg <= dl_in_vec;
            end
        end
    end
    
    // find_df_deadlock to report the deadlock
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            find_df_deadlock <= 1'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED && dl_detect_reg == dl_done_reg) begin
                find_df_deadlock <= 1'b1;
            end
            else if (CS_fsm == ST_IDLE) begin
                find_df_deadlock <= 1'b0;
            end
        end
    end
    
    // get the first valid proc index in dl vector
    function integer proc_index(input [PROC_NUM - 1:0] dl_vec);
        begin
            proc_index = 0;
            for (i = 0; i < PROC_NUM; i = i + 1) begin
                if (dl_vec[i]) begin
                    proc_index = i;
                end
            end
        end
    endfunction

    // get the proc path based on dl vector
    function [304:0] proc_path(input [PROC_NUM - 1:0] dl_vec);
        integer index;
        begin
            index = proc_index(dl_vec);
            case (index)
                0 : begin
                    proc_path = "top.entry_proc_U0";
                end
                1 : begin
                    proc_path = "top.Block_entry3_proc_U0";
                end
                2 : begin
                    proc_path = "top.ConvertBias_BN_U0";
                end
                3 : begin
                    proc_path = "top.ConvertInputToStream_U0";
                end
                4 : begin
                    proc_path = "top.Padding_U0";
                end
                5 : begin
                    proc_path = "top.Sliding_U0";
                end
                6 : begin
                    proc_path = "top.ConvertInputToArray_U0";
                end
                7 : begin
                    proc_path = "top.ConvertWeightToStream_U0";
                end
                8 : begin
                    proc_path = "top.ConvWeightToArray_U0";
                end
                9 : begin
                    proc_path = "top.MMWeightToArray_U0";
                end
                10 : begin
                    proc_path = "top.MuxWeightStream_U0";
                end
                11 : begin
                    proc_path = "top.Compute_U0";
                end
                12 : begin
                    proc_path = "top.ConvertToOutStream_U0";
                end
                13 : begin
                    proc_path = "top.ConvToOutStream_U0";
                end
                14 : begin
                    proc_path = "top.ConvBias_U0";
                end
                15 : begin
                    proc_path = "top.ConvBN_U0";
                end
                16 : begin
                    proc_path = "top.ResOutput_U0";
                end
                default : begin
                    proc_path = "unknown";
                end
            endcase
        end
    endfunction

    // print the headlines of deadlock detection
    task print_dl_head;
        begin
            $display("\n//////////////////////////////////////////////////////////////////////////////");
            $display("// ERROR!!! DEADLOCK DETECTED at %0t ns! SIMULATION WILL BE STOPPED! //", $time);
            $display("//////////////////////////////////////////////////////////////////////////////");
            fp = $fopen("deadlock_db.dat", "w");
        end
    endtask

    // print the start of a cycle
    task print_cycle_start(input reg [304:0] proc_path, input integer cycle_id);
        begin
            $display("/////////////////////////");
            $display("// Dependence cycle %0d:", cycle_id);
            $display("// (1): Process: %0s", proc_path);
            $fdisplay(fp, "Dependence_Cycle_ID %0d", cycle_id);
            $fdisplay(fp, "Dependence_Process_ID 1");
            $fdisplay(fp, "Dependence_Process_path %0s", proc_path);
        end
    endtask

    // print the end of deadlock detection
    task print_dl_end(input integer num, input integer record_time);
        begin
            $display("////////////////////////////////////////////////////////////////////////");
            $display("// Totally %0d cycles detected!", num);
            $display("////////////////////////////////////////////////////////////////////////");
            $fdisplay(fp, "Dependence_Cycle_Number %0d", num);
            $fclose(fp);
        end
    endtask

    // print one proc component in the cycle
    task print_cycle_proc_comp(input reg [304:0] proc_path, input integer cycle_comp_id);
        begin
            $display("// (%0d): Process: %0s", cycle_comp_id, proc_path);
            $fdisplay(fp, "Dependence_Process_ID %0d", cycle_comp_id);
            $fdisplay(fp, "Dependence_Process_path %0s", proc_path);
        end
    endtask

    // print one channel component in the cycle
    task print_cycle_chan_comp(input [PROC_NUM - 1:0] dl_vec1, input [PROC_NUM - 1:0] dl_vec2);
        reg [376:0] chan_path;
        integer index1;
        integer index2;
        begin
            index1 = proc_index(dl_vec1);
            index2 = proc_index(dl_vec2);
            case (index1)
                0 : begin
                    case(index2)
                    16: begin
                        if (~AESL_inst_top.entry_proc_U0.Output_r_c_blk_n) begin
                            if (~AESL_inst_top.Output_r_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Output_r_c_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Output_r_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Output_r_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Output_r_c_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Output_r_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.start_for_ResOutput_U0_U.if_full_n & AESL_inst_top.entry_proc_U0.ap_start & ~AESL_inst_top.entry_proc_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~AESL_inst_top.start_for_ResOutput_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'top.start_for_ResOutput_U0_U' read by process 'top.ResOutput_U0',");
                        end
                    end
                    5: begin
                        if (~AESL_inst_top.entry_proc_U0.K_c58_blk_n) begin
                            if (~AESL_inst_top.K_c58_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.K_c58_U' written by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.K_c58_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.K_c58_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.K_c58_U' read by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.K_c58_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.entry_proc_U0.S_c61_blk_n) begin
                            if (~AESL_inst_top.S_c61_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.S_c61_U' written by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.S_c61_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.S_c61_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.S_c61_U' read by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.S_c61_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.start_for_Sliding_U0_U.if_full_n & AESL_inst_top.entry_proc_U0.ap_start & ~AESL_inst_top.entry_proc_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~AESL_inst_top.start_for_Sliding_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'top.start_for_Sliding_U0_U' read by process 'top.Sliding_U0',");
                        end
                    end
                    4: begin
                        if (~AESL_inst_top.entry_proc_U0.P_c60_blk_n) begin
                            if (~AESL_inst_top.P_c60_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.P_c60_U' written by process 'top.Padding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.P_c60_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.P_c60_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.P_c60_U' read by process 'top.Padding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.P_c60_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.start_for_Padding_U0_U.if_full_n & AESL_inst_top.entry_proc_U0.ap_start & ~AESL_inst_top.entry_proc_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~AESL_inst_top.start_for_Padding_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'top.start_for_Padding_U0_U' read by process 'top.Padding_U0',");
                        end
                    end
                    1: begin
                        if (AESL_inst_top.ap_sync_entry_proc_U0_ap_ready & AESL_inst_top.entry_proc_U0.ap_idle & ~AESL_inst_top.ap_sync_Block_entry3_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'top.Block_entry3_proc_U0'");
                        end
                    end
                    2: begin
                        if (AESL_inst_top.ap_sync_entry_proc_U0_ap_ready & AESL_inst_top.entry_proc_U0.ap_idle & ~AESL_inst_top.ap_sync_ConvertBias_BN_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'top.ConvertBias_BN_U0'");
                        end
                    end
                    3: begin
                        if (AESL_inst_top.ap_sync_entry_proc_U0_ap_ready & AESL_inst_top.entry_proc_U0.ap_idle & ~AESL_inst_top.ap_sync_ConvertInputToStream_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'top.ConvertInputToStream_U0'");
                        end
                    end
                    7: begin
                        if (AESL_inst_top.ap_sync_entry_proc_U0_ap_ready & AESL_inst_top.entry_proc_U0.ap_idle & ~AESL_inst_top.ap_sync_ConvertWeightToStream_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'top.ConvertWeightToStream_U0'");
                        end
                    end
                    endcase
                end
                1 : begin
                    case(index2)
                    0: begin
                        if (AESL_inst_top.ap_sync_Block_entry3_proc_U0_ap_ready & AESL_inst_top.Block_entry3_proc_U0.ap_idle & ~AESL_inst_top.ap_sync_entry_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'top.entry_proc_U0'");
                        end
                    end
                    2: begin
                        if (AESL_inst_top.ap_sync_Block_entry3_proc_U0_ap_ready & AESL_inst_top.Block_entry3_proc_U0.ap_idle & ~AESL_inst_top.ap_sync_ConvertBias_BN_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'top.ConvertBias_BN_U0'");
                        end
                    end
                    3: begin
                        if (AESL_inst_top.ap_sync_Block_entry3_proc_U0_ap_ready & AESL_inst_top.Block_entry3_proc_U0.ap_idle & ~AESL_inst_top.ap_sync_ConvertInputToStream_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'top.ConvertInputToStream_U0'");
                        end
                    end
                    7: begin
                        if (AESL_inst_top.ap_sync_Block_entry3_proc_U0_ap_ready & AESL_inst_top.Block_entry3_proc_U0.ap_idle & ~AESL_inst_top.ap_sync_ConvertWeightToStream_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'top.ConvertWeightToStream_U0'");
                        end
                    end
                    endcase
                end
                2 : begin
                    case(index2)
                    15: begin
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_0_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_1_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_1_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_1_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_2_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_2_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_2_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_3_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_3_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_3_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_4_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_4_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_4_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_5_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_5_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_5_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_6_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_6_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_6_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_7_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_7_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_7_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_8_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_8_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_8_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_9_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_9_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_9_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_10_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_10_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_10_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_11_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_11_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_11_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_12_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_12_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_12_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_13_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_13_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_13_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_14_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_14_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_14_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_15_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_15_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_15_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_16_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_16_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_16_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_17_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_17_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_17_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_18_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_18_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_18_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_19_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_19_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_19_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_20_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_20_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_20_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_21_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_21_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_21_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_22_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_22_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_22_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_23_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_23_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_23_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_24_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_24_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_24_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_25_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_25_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_25_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_26_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_26_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_26_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_27_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_27_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_27_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_28_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_28_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_28_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_29_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_29_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_29_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_30_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_30_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_30_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_31_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_31_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_31_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_32_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_32_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_32_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_33_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_33_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_33_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_34_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_34_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_34_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_35_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_35_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_35_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_36_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_36_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_36_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_37_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_37_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_37_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_38_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_38_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_38_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_39_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_39_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_39_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_40_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_40_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_40_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_40_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_40_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_40_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_40_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_41_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_41_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_41_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_41_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_41_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_41_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_41_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_42_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_42_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_42_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_42_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_42_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_42_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_42_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_43_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_43_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_43_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_43_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_43_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_43_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_43_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_44_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_44_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_44_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_44_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_44_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_44_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_44_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_45_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_45_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_45_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_45_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_45_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_45_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_45_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_46_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_46_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_46_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_46_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_46_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_46_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_46_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_47_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_47_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_47_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_47_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_47_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_47_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_47_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_48_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_48_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_48_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_48_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_48_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_48_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_48_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_49_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_49_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_49_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_49_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_49_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_49_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_49_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_50_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_50_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_50_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_50_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_50_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_50_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_50_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_51_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_51_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_51_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_51_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_51_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_51_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_51_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_52_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_52_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_52_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_52_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_52_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_52_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_52_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_53_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_53_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_53_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_53_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_53_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_53_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_53_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_54_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_54_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_54_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_54_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_54_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_54_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_54_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_55_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_55_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_55_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_55_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_55_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_55_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_55_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_56_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_56_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_56_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_56_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_56_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_56_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_56_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_57_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_57_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_57_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_57_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_57_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_57_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_57_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_58_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_58_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_58_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_58_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_58_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_58_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_58_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_59_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_59_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_59_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_59_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_59_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_59_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_59_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_60_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_60_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_60_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_60_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_60_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_60_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_60_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_61_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_61_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_61_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_61_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_61_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_61_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_61_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_62_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_62_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_62_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_62_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_62_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_62_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_62_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_63_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_63_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_63_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_63_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_63_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_63_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_63_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_64_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_64_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_64_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_64_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_64_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_64_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_64_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_65_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_65_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_65_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_65_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_65_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_65_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_65_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_66_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_66_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_66_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_66_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_66_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_66_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_66_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_67_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_67_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_67_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_67_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_67_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_67_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_67_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_68_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_68_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_68_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_68_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_68_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_68_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_68_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_69_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_69_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_69_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_69_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_69_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_69_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_69_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_70_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_70_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_70_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_70_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_70_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_70_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_70_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_71_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_71_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_71_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_71_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_71_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_71_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_71_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_72_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_72_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_72_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_72_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_72_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_72_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_72_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_73_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_73_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_73_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_73_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_73_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_73_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_73_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_74_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_74_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_74_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_74_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_74_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_74_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_74_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_75_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_75_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_75_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_75_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_75_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_75_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_75_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_76_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_76_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_76_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_76_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_76_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_76_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_76_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_77_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_77_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_77_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_77_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_77_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_77_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_77_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_78_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_78_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_78_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_78_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_78_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_78_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_78_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_79_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_79_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_79_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_79_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_79_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_79_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_79_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_80_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_80_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_80_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_80_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_80_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_80_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_80_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_81_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_81_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_81_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_81_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_81_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_81_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_81_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_82_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_82_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_82_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_82_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_82_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_82_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_82_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_83_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_83_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_83_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_83_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_83_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_83_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_83_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_84_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_84_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_84_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_84_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_84_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_84_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_84_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_85_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_85_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_85_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_85_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_85_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_85_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_85_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_86_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_86_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_86_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_86_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_86_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_86_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_86_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_87_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_87_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_87_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_87_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_87_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_87_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_87_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_88_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_88_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_88_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_88_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_88_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_88_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_88_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_89_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_89_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_89_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_89_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_89_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_89_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_89_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_90_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_90_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_90_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_90_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_90_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_90_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_90_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_91_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_91_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_91_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_91_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_91_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_91_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_91_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_92_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_92_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_92_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_92_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_92_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_92_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_92_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_93_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_93_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_93_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_93_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_93_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_93_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_93_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_94_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_94_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_94_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_94_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_94_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_94_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_94_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_95_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_95_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_95_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_95_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_95_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_95_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_95_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_96_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_96_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_96_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_96_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_96_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_96_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_96_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_97_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_97_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_97_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_97_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_97_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_97_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_97_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_98_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_98_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_98_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_98_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_98_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_98_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_98_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_99_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_99_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_99_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_99_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_99_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_99_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_99_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_100_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_100_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_100_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_100_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_100_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_100_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_100_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_101_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_101_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_101_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_101_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_101_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_101_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_101_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_102_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_102_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_102_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_102_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_102_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_102_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_102_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_103_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_103_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_103_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_103_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_103_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_103_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_103_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_104_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_104_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_104_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_104_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_104_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_104_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_104_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_105_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_105_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_105_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_105_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_105_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_105_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_105_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_106_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_106_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_106_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_106_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_106_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_106_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_106_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_107_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_107_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_107_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_107_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_107_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_107_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_107_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_108_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_108_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_108_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_108_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_108_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_108_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_108_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_109_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_109_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_109_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_109_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_109_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_109_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_109_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_110_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_110_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_110_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_110_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_110_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_110_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_110_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_111_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_111_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_111_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_111_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_111_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_111_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_111_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_112_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_112_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_112_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_112_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_112_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_112_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_112_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_113_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_113_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_113_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_113_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_113_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_113_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_113_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_114_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_114_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_114_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_114_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_114_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_114_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_114_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_115_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_115_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_115_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_115_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_115_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_115_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_115_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_116_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_116_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_116_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_116_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_116_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_116_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_116_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_117_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_117_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_117_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_117_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_117_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_117_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_117_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_118_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_118_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_118_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_118_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_118_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_118_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_118_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_119_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_119_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_119_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_119_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_119_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_119_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_119_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_120_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_120_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_120_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_120_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_120_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_120_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_120_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_121_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_121_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_121_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_121_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_121_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_121_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_121_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_122_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_122_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_122_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_122_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_122_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_122_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_122_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_123_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_123_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_123_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_123_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_123_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_123_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_123_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_124_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_124_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_124_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_124_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_124_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_124_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_124_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_125_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_125_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_125_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_125_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_125_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_125_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_125_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_126_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_126_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_126_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_126_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_126_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_126_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_126_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_norm_127_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_127_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_127_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_127_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_127_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_127_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_127_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.start_for_ConvBN_U0_U.if_full_n & AESL_inst_top.ConvertBias_BN_U0.ap_start & ~AESL_inst_top.ConvertBias_BN_U0.real_start & (trans_in_cnt_3 == trans_out_cnt_3) & ~AESL_inst_top.start_for_ConvBN_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'top.start_for_ConvBN_U0_U' read by process 'top.ConvBN_U0',");
                        end
                    end
                    14: begin
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_0_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_1_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_1_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_1_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_2_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_2_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_2_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_3_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_3_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_3_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_4_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_4_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_4_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_5_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_5_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_5_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_6_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_6_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_6_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_7_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_7_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_7_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_8_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_8_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_8_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_9_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_9_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_9_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_10_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_10_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_10_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_11_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_11_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_11_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_12_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_12_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_12_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_13_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_13_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_13_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_14_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_14_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_14_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_15_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_15_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_15_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_16_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_16_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_16_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_17_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_17_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_17_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_18_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_18_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_18_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_19_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_19_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_19_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_20_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_20_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_20_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_21_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_21_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_21_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_22_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_22_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_22_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_23_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_23_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_23_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_24_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_24_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_24_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_25_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_25_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_25_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_26_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_26_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_26_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_27_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_27_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_27_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_28_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_28_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_28_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_29_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_29_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_29_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_30_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_30_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_30_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_31_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_31_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_31_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_32_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_32_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_32_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_33_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_33_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_33_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_34_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_34_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_34_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_35_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_35_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_35_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_36_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_36_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_36_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_37_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_37_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_37_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_38_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_38_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_38_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_39_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_39_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_39_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_40_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_40_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_40_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_40_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_40_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_40_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_40_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_41_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_41_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_41_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_41_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_41_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_41_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_41_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_42_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_42_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_42_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_42_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_42_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_42_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_42_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_43_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_43_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_43_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_43_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_43_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_43_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_43_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_44_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_44_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_44_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_44_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_44_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_44_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_44_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_45_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_45_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_45_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_45_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_45_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_45_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_45_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_46_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_46_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_46_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_46_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_46_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_46_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_46_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_47_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_47_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_47_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_47_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_47_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_47_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_47_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_48_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_48_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_48_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_48_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_48_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_48_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_48_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_49_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_49_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_49_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_49_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_49_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_49_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_49_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_50_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_50_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_50_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_50_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_50_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_50_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_50_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_51_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_51_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_51_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_51_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_51_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_51_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_51_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_52_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_52_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_52_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_52_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_52_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_52_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_52_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_53_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_53_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_53_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_53_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_53_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_53_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_53_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_54_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_54_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_54_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_54_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_54_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_54_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_54_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_55_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_55_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_55_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_55_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_55_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_55_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_55_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_56_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_56_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_56_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_56_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_56_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_56_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_56_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_57_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_57_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_57_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_57_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_57_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_57_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_57_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_58_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_58_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_58_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_58_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_58_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_58_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_58_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_59_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_59_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_59_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_59_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_59_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_59_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_59_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_60_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_60_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_60_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_60_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_60_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_60_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_60_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_61_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_61_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_61_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_61_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_61_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_61_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_61_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_62_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_62_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_62_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_62_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_62_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_62_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_62_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_63_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_63_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_63_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_63_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_63_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_63_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_63_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_64_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_64_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_64_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_64_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_64_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_64_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_64_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_65_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_65_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_65_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_65_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_65_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_65_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_65_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_66_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_66_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_66_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_66_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_66_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_66_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_66_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_67_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_67_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_67_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_67_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_67_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_67_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_67_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_68_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_68_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_68_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_68_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_68_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_68_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_68_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_69_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_69_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_69_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_69_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_69_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_69_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_69_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_70_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_70_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_70_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_70_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_70_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_70_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_70_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_71_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_71_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_71_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_71_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_71_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_71_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_71_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_72_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_72_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_72_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_72_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_72_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_72_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_72_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_73_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_73_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_73_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_73_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_73_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_73_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_73_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_74_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_74_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_74_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_74_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_74_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_74_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_74_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_75_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_75_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_75_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_75_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_75_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_75_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_75_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_76_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_76_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_76_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_76_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_76_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_76_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_76_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_77_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_77_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_77_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_77_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_77_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_77_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_77_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_78_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_78_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_78_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_78_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_78_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_78_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_78_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_79_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_79_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_79_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_79_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_79_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_79_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_79_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_80_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_80_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_80_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_80_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_80_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_80_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_80_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_81_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_81_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_81_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_81_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_81_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_81_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_81_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_82_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_82_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_82_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_82_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_82_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_82_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_82_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_83_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_83_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_83_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_83_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_83_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_83_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_83_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_84_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_84_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_84_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_84_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_84_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_84_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_84_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_85_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_85_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_85_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_85_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_85_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_85_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_85_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_86_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_86_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_86_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_86_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_86_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_86_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_86_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_87_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_87_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_87_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_87_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_87_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_87_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_87_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_88_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_88_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_88_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_88_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_88_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_88_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_88_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_89_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_89_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_89_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_89_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_89_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_89_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_89_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_90_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_90_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_90_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_90_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_90_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_90_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_90_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_91_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_91_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_91_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_91_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_91_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_91_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_91_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_92_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_92_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_92_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_92_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_92_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_92_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_92_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_93_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_93_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_93_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_93_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_93_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_93_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_93_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_94_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_94_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_94_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_94_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_94_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_94_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_94_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_95_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_95_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_95_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_95_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_95_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_95_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_95_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_96_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_96_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_96_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_96_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_96_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_96_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_96_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_97_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_97_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_97_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_97_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_97_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_97_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_97_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_98_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_98_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_98_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_98_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_98_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_98_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_98_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_99_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_99_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_99_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_99_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_99_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_99_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_99_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_100_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_100_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_100_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_100_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_100_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_100_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_100_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_101_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_101_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_101_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_101_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_101_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_101_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_101_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_102_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_102_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_102_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_102_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_102_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_102_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_102_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_103_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_103_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_103_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_103_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_103_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_103_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_103_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_104_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_104_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_104_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_104_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_104_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_104_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_104_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_105_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_105_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_105_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_105_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_105_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_105_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_105_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_106_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_106_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_106_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_106_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_106_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_106_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_106_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_107_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_107_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_107_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_107_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_107_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_107_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_107_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_108_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_108_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_108_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_108_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_108_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_108_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_108_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_109_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_109_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_109_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_109_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_109_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_109_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_109_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_110_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_110_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_110_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_110_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_110_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_110_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_110_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_111_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_111_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_111_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_111_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_111_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_111_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_111_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_112_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_112_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_112_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_112_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_112_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_112_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_112_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_113_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_113_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_113_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_113_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_113_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_113_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_113_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_114_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_114_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_114_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_114_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_114_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_114_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_114_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_115_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_115_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_115_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_115_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_115_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_115_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_115_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_116_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_116_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_116_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_116_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_116_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_116_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_116_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_117_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_117_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_117_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_117_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_117_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_117_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_117_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_118_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_118_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_118_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_118_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_118_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_118_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_118_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_119_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_119_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_119_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_119_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_119_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_119_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_119_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_120_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_120_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_120_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_120_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_120_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_120_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_120_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_121_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_121_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_121_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_121_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_121_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_121_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_121_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_122_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_122_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_122_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_122_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_122_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_122_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_122_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_123_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_123_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_123_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_123_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_123_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_123_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_123_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_124_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_124_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_124_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_124_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_124_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_124_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_124_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_125_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_125_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_125_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_125_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_125_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_125_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_125_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_126_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_126_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_126_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_126_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_126_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_126_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_126_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertBias_BN_U0.grp_ConvertBias_BN_Pipeline_VITIS_LOOP_7_1_fu_566.fifo_bias_127_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_127_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_127_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_127_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_127_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_127_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_127_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.start_for_ConvBias_U0_U.if_full_n & AESL_inst_top.ConvertBias_BN_U0.ap_start & ~AESL_inst_top.ConvertBias_BN_U0.real_start & (trans_in_cnt_3 == trans_out_cnt_3) & ~AESL_inst_top.start_for_ConvBias_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'top.start_for_ConvBias_U0_U' read by process 'top.ConvBias_U0',");
                        end
                    end
                    0: begin
                        if (AESL_inst_top.ap_sync_ConvertBias_BN_U0_ap_ready & AESL_inst_top.ConvertBias_BN_U0.ap_idle & ~AESL_inst_top.ap_sync_entry_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'top.entry_proc_U0'");
                        end
                    end
                    1: begin
                        if (AESL_inst_top.ap_sync_ConvertBias_BN_U0_ap_ready & AESL_inst_top.ConvertBias_BN_U0.ap_idle & ~AESL_inst_top.ap_sync_Block_entry3_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'top.Block_entry3_proc_U0'");
                        end
                    end
                    3: begin
                        if (AESL_inst_top.ap_sync_ConvertBias_BN_U0_ap_ready & AESL_inst_top.ConvertBias_BN_U0.ap_idle & ~AESL_inst_top.ap_sync_ConvertInputToStream_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'top.ConvertInputToStream_U0'");
                        end
                    end
                    7: begin
                        if (AESL_inst_top.ap_sync_ConvertBias_BN_U0_ap_ready & AESL_inst_top.ConvertBias_BN_U0.ap_idle & ~AESL_inst_top.ap_sync_ConvertWeightToStream_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'top.ConvertWeightToStream_U0'");
                        end
                    end
                    endcase
                end
                3 : begin
                    case(index2)
                    4: begin
                        if (~AESL_inst_top.ConvertInputToStream_U0.grp_ConvertInputToStream_Pipeline_VITIS_LOOP_19_1_VITIS_LOOP_22_2_VITIS_LOOP_25_3_VI_fu_166.conv_a_blk_n) begin
                            if (~AESL_inst_top.conv_a_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.conv_a_U' written by process 'top.Padding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.conv_a_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.conv_a_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.conv_a_U' read by process 'top.Padding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.conv_a_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertInputToStream_U0.R_c46_blk_n) begin
                            if (~AESL_inst_top.R_c46_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.R_c46_U' written by process 'top.Padding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.R_c46_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.R_c46_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.R_c46_U' read by process 'top.Padding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.R_c46_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertInputToStream_U0.C_c48_blk_n) begin
                            if (~AESL_inst_top.C_c48_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.C_c48_U' written by process 'top.Padding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.C_c48_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.C_c48_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.C_c48_U' read by process 'top.Padding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.C_c48_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertInputToStream_U0.N_c51_blk_n) begin
                            if (~AESL_inst_top.N_c51_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.N_c51_U' written by process 'top.Padding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.N_c51_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.N_c51_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.N_c51_U' read by process 'top.Padding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.N_c51_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertInputToStream_U0.M_c56_blk_n) begin
                            if (~AESL_inst_top.M_c56_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.M_c56_U' written by process 'top.Padding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.M_c56_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.M_c56_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.M_c56_U' read by process 'top.Padding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.M_c56_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertInputToStream_U0.mode_c72_blk_n) begin
                            if (~AESL_inst_top.mode_c72_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.mode_c72_U' written by process 'top.Padding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c72_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.mode_c72_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.mode_c72_U' read by process 'top.Padding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c72_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    6: begin
                        if (~AESL_inst_top.ConvertInputToStream_U0.grp_ConvertInputToStream_Pipeline_VITIS_LOOP_40_5_VITIS_LOOP_43_6_VITIS_LOOP_46_7_fu_154.mm_a_blk_n) begin
                            if (~AESL_inst_top.mm_a_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.mm_a_U' written by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mm_a_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.mm_a_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.mm_a_U' read by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mm_a_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    0: begin
                        if (AESL_inst_top.ap_sync_ConvertInputToStream_U0_ap_ready & AESL_inst_top.ConvertInputToStream_U0.ap_idle & ~AESL_inst_top.ap_sync_entry_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'top.entry_proc_U0'");
                        end
                    end
                    1: begin
                        if (AESL_inst_top.ap_sync_ConvertInputToStream_U0_ap_ready & AESL_inst_top.ConvertInputToStream_U0.ap_idle & ~AESL_inst_top.ap_sync_Block_entry3_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'top.Block_entry3_proc_U0'");
                        end
                    end
                    2: begin
                        if (AESL_inst_top.ap_sync_ConvertInputToStream_U0_ap_ready & AESL_inst_top.ConvertInputToStream_U0.ap_idle & ~AESL_inst_top.ap_sync_ConvertBias_BN_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'top.ConvertBias_BN_U0'");
                        end
                    end
                    7: begin
                        if (AESL_inst_top.ap_sync_ConvertInputToStream_U0_ap_ready & AESL_inst_top.ConvertInputToStream_U0.ap_idle & ~AESL_inst_top.ap_sync_ConvertWeightToStream_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'top.ConvertWeightToStream_U0'");
                        end
                    end
                    endcase
                end
                4 : begin
                    case(index2)
                    3: begin
                        if (~AESL_inst_top.Padding_U0.grp_Padding_Pipeline_VITIS_LOOP_62_1_VITIS_LOOP_65_2_VITIS_LOOP_68_3_VITIS_LOOP_71_4_fu_152.conv_a_blk_n) begin
                            if (~AESL_inst_top.conv_a_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.conv_a_U' written by process 'top.ConvertInputToStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.conv_a_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.conv_a_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.conv_a_U' read by process 'top.ConvertInputToStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.conv_a_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Padding_U0.R_blk_n) begin
                            if (~AESL_inst_top.R_c46_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.R_c46_U' written by process 'top.ConvertInputToStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.R_c46_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.R_c46_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.R_c46_U' read by process 'top.ConvertInputToStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.R_c46_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Padding_U0.C_blk_n) begin
                            if (~AESL_inst_top.C_c48_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.C_c48_U' written by process 'top.ConvertInputToStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.C_c48_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.C_c48_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.C_c48_U' read by process 'top.ConvertInputToStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.C_c48_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Padding_U0.N_blk_n) begin
                            if (~AESL_inst_top.N_c51_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.N_c51_U' written by process 'top.ConvertInputToStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.N_c51_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.N_c51_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.N_c51_U' read by process 'top.ConvertInputToStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.N_c51_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Padding_U0.M_blk_n) begin
                            if (~AESL_inst_top.M_c56_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.M_c56_U' written by process 'top.ConvertInputToStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.M_c56_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.M_c56_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.M_c56_U' read by process 'top.ConvertInputToStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.M_c56_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Padding_U0.mode_blk_n) begin
                            if (~AESL_inst_top.mode_c72_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.mode_c72_U' written by process 'top.ConvertInputToStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c72_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.mode_c72_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.mode_c72_U' read by process 'top.ConvertInputToStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c72_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    5: begin
                        if (~AESL_inst_top.Padding_U0.grp_Padding_Pipeline_VITIS_LOOP_62_1_VITIS_LOOP_65_2_VITIS_LOOP_68_3_VITIS_LOOP_71_4_fu_152.conv3_samepad_blk_n) begin
                            if (~AESL_inst_top.conv3_samepad_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.conv3_samepad_U' written by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.conv3_samepad_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.conv3_samepad_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.conv3_samepad_U' read by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.conv3_samepad_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Padding_U0.R_c45_blk_n) begin
                            if (~AESL_inst_top.R_c45_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.R_c45_U' written by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.R_c45_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.R_c45_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.R_c45_U' read by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.R_c45_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Padding_U0.C_c47_blk_n) begin
                            if (~AESL_inst_top.C_c47_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.C_c47_U' written by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.C_c47_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.C_c47_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.C_c47_U' read by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.C_c47_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Padding_U0.N_c50_blk_n) begin
                            if (~AESL_inst_top.N_c50_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.N_c50_U' written by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.N_c50_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.N_c50_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.N_c50_U' read by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.N_c50_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Padding_U0.M_c55_blk_n) begin
                            if (~AESL_inst_top.M_c55_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.M_c55_U' written by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.M_c55_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.M_c55_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.M_c55_U' read by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.M_c55_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Padding_U0.P_c59_blk_n) begin
                            if (~AESL_inst_top.P_c59_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.P_c59_U' written by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.P_c59_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.P_c59_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.P_c59_U' read by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.P_c59_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Padding_U0.mode_c71_blk_n) begin
                            if (~AESL_inst_top.mode_c71_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.mode_c71_U' written by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c71_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.mode_c71_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.mode_c71_U' read by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c71_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    0: begin
                        if (~AESL_inst_top.Padding_U0.P_blk_n) begin
                            if (~AESL_inst_top.P_c60_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.P_c60_U' written by process 'top.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.P_c60_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.P_c60_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.P_c60_U' read by process 'top.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.P_c60_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.start_for_Padding_U0_U.if_empty_n & AESL_inst_top.Padding_U0.ap_idle & ~AESL_inst_top.start_for_Padding_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'top.start_for_Padding_U0_U' written by process 'top.entry_proc_U0',");
                        end
                    end
                    endcase
                end
                5 : begin
                    case(index2)
                    4: begin
                        if (~AESL_inst_top.Sliding_U0.grp_Sliding_Pipeline_VITIS_LOOP_114_1_VITIS_LOOP_117_2_fu_192.conv3_samepad_blk_n) begin
                            if (~AESL_inst_top.conv3_samepad_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.conv3_samepad_U' written by process 'top.Padding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.conv3_samepad_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.conv3_samepad_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.conv3_samepad_U' read by process 'top.Padding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.conv3_samepad_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Sliding_U0.R_blk_n) begin
                            if (~AESL_inst_top.R_c45_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.R_c45_U' written by process 'top.Padding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.R_c45_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.R_c45_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.R_c45_U' read by process 'top.Padding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.R_c45_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Sliding_U0.C_blk_n) begin
                            if (~AESL_inst_top.C_c47_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.C_c47_U' written by process 'top.Padding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.C_c47_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.C_c47_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.C_c47_U' read by process 'top.Padding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.C_c47_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Sliding_U0.N_blk_n) begin
                            if (~AESL_inst_top.N_c50_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.N_c50_U' written by process 'top.Padding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.N_c50_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.N_c50_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.N_c50_U' read by process 'top.Padding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.N_c50_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Sliding_U0.M_blk_n) begin
                            if (~AESL_inst_top.M_c55_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.M_c55_U' written by process 'top.Padding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.M_c55_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.M_c55_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.M_c55_U' read by process 'top.Padding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.M_c55_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Sliding_U0.P_blk_n) begin
                            if (~AESL_inst_top.P_c59_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.P_c59_U' written by process 'top.Padding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.P_c59_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.P_c59_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.P_c59_U' read by process 'top.Padding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.P_c59_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Sliding_U0.mode_blk_n) begin
                            if (~AESL_inst_top.mode_c71_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.mode_c71_U' written by process 'top.Padding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c71_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.mode_c71_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.mode_c71_U' read by process 'top.Padding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c71_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    6: begin
                        if (~AESL_inst_top.Sliding_U0.grp_Sliding_Pipeline_VITIS_LOOP_114_1_VITIS_LOOP_117_2_fu_192.conv3_sild_blk_n) begin
                            if (~AESL_inst_top.conv3_sild_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.conv3_sild_U' written by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.conv3_sild_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.conv3_sild_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.conv3_sild_U' read by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.conv3_sild_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Sliding_U0.mode_c70_blk_n) begin
                            if (~AESL_inst_top.mode_c70_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.mode_c70_U' written by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c70_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.mode_c70_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.mode_c70_U' read by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c70_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    0: begin
                        if (~AESL_inst_top.Sliding_U0.K_blk_n) begin
                            if (~AESL_inst_top.K_c58_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.K_c58_U' written by process 'top.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.K_c58_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.K_c58_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.K_c58_U' read by process 'top.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.K_c58_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Sliding_U0.S_blk_n) begin
                            if (~AESL_inst_top.S_c61_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.S_c61_U' written by process 'top.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.S_c61_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.S_c61_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.S_c61_U' read by process 'top.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.S_c61_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.start_for_Sliding_U0_U.if_empty_n & AESL_inst_top.Sliding_U0.ap_idle & ~AESL_inst_top.start_for_Sliding_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'top.start_for_Sliding_U0_U' written by process 'top.entry_proc_U0',");
                        end
                    end
                    12: begin
                        if (~AESL_inst_top.Sliding_U0.R_c44_blk_n) begin
                            if (~AESL_inst_top.R_c44_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.R_c44_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.R_c44_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.R_c44_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.R_c44_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.R_c44_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Sliding_U0.N_c49_blk_n) begin
                            if (~AESL_inst_top.N_c49_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.N_c49_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.N_c49_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.N_c49_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.N_c49_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.N_c49_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.start_for_ConvertToOutStream_U0_U.if_full_n & AESL_inst_top.Sliding_U0.ap_start & ~AESL_inst_top.Sliding_U0.real_start & (trans_in_cnt_2 == trans_out_cnt_2) & ~AESL_inst_top.start_for_ConvertToOutStream_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'top.start_for_ConvertToOutStream_U0_U' read by process 'top.ConvertToOutStream_U0',");
                        end
                    end
                    16: begin
                        if (~AESL_inst_top.Sliding_U0.C_c_blk_n) begin
                            if (~AESL_inst_top.C_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.C_c_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.C_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.C_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.C_c_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.C_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Sliding_U0.P_c_blk_n) begin
                            if (~AESL_inst_top.P_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.P_c_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.P_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.P_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.P_c_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.P_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Sliding_U0.S_c_blk_n) begin
                            if (~AESL_inst_top.S_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.S_c_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.S_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.S_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.S_c_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.S_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    13: begin
                        if (~AESL_inst_top.Sliding_U0.M_c54_blk_n) begin
                            if (~AESL_inst_top.M_c54_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.M_c54_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.M_c54_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.M_c54_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.M_c54_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.M_c54_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Sliding_U0.K_c57_blk_n) begin
                            if (~AESL_inst_top.K_c57_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.K_c57_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.K_c57_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.K_c57_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.K_c57_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.K_c57_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                6 : begin
                    case(index2)
                    5: begin
                        if (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.conv3_sild_blk_n) begin
                            if (~AESL_inst_top.conv3_sild_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.conv3_sild_U' written by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.conv3_sild_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.conv3_sild_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.conv3_sild_U' read by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.conv3_sild_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertInputToArray_U0.mode_blk_n) begin
                            if (~AESL_inst_top.mode_c70_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.mode_c70_U' written by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c70_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.mode_c70_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.mode_c70_U' read by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c70_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    3: begin
                        if (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.mm_a_blk_n) begin
                            if (~AESL_inst_top.mm_a_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.mm_a_U' written by process 'top.ConvertInputToStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mm_a_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.mm_a_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.mm_a_U' read by process 'top.ConvertInputToStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mm_a_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    11: begin
                        if (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.fifo_SA_A_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_A_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_A_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_A_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_A_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.fifo_SA_A_1_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_A_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_A_1_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_A_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_A_1_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.fifo_SA_A_2_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_A_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_A_2_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_A_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_A_2_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.fifo_SA_A_3_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_A_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_A_3_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_A_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_A_3_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.fifo_SA_A_4_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_A_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_A_4_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_A_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_A_4_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.fifo_SA_A_5_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_A_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_A_5_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_A_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_A_5_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.fifo_SA_A_6_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_A_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_A_6_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_A_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_A_6_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.fifo_SA_A_7_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_A_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_A_7_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_A_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_A_7_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.fifo_SA_A_8_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_A_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_A_8_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_A_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_A_8_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.fifo_SA_A_9_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_A_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_A_9_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_A_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_A_9_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.fifo_SA_A_10_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_A_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_A_10_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_A_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_A_10_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.fifo_SA_A_11_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_A_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_A_11_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_A_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_A_11_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.fifo_SA_A_12_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_A_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_A_12_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_A_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_A_12_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.fifo_SA_A_13_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_A_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_A_13_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_A_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_A_13_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.fifo_SA_A_14_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_A_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_A_14_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_A_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_A_14_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertInputToArray_U0.grp_ConvertInputToArray_Pipeline_VITIS_LOOP_201_1_fu_104.fifo_SA_A_15_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_A_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_A_15_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_A_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_A_15_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertInputToArray_U0.num_a_sa_2_loc_c42_blk_n) begin
                            if (~AESL_inst_top.num_a_sa_2_loc_c42_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.num_a_sa_2_loc_c42_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.num_a_sa_2_loc_c42_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.num_a_sa_2_loc_c42_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.num_a_sa_2_loc_c42_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.num_a_sa_2_loc_c42_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertInputToArray_U0.mode_c66_blk_n) begin
                            if (~AESL_inst_top.mode_c66_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.mode_c66_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c66_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.mode_c66_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.mode_c66_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c66_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    1: begin
                        if (~AESL_inst_top.num_a_sa_2_loc_c43_channel_U.if_empty_n & AESL_inst_top.ConvertInputToArray_U0.ap_idle & ~AESL_inst_top.num_a_sa_2_loc_c43_channel_U.if_write) begin
                            if (~AESL_inst_top.num_a_sa_2_loc_c43_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.num_a_sa_2_loc_c43_channel_U' written by process 'top.Block_entry3_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.num_a_sa_2_loc_c43_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.num_a_sa_2_loc_c43_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.num_a_sa_2_loc_c43_channel_U' read by process 'top.Block_entry3_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.num_a_sa_2_loc_c43_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                7 : begin
                    case(index2)
                    8: begin
                        if (~AESL_inst_top.ConvertWeightToStream_U0.grp_ConvertWeightToStream_Pipeline_VITIS_LOOP_229_1_VITIS_LOOP_232_2_VITIS_LOOP_234_s_fu_180.fifo_conv_w_0_blk_n) begin
                            if (~AESL_inst_top.fifo_conv_w_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_conv_w_U' written by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_conv_w_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_conv_w_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_conv_w_U' read by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_conv_w_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertWeightToStream_U0.grp_ConvertWeightToStream_Pipeline_VITIS_LOOP_229_1_VITIS_LOOP_232_2_VITIS_LOOP_234_s_fu_180.fifo_conv_w_1_blk_n) begin
                            if (~AESL_inst_top.fifo_conv_w_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_conv_w_1_U' written by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_conv_w_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_conv_w_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_conv_w_1_U' read by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_conv_w_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertWeightToStream_U0.grp_ConvertWeightToStream_Pipeline_VITIS_LOOP_229_1_VITIS_LOOP_232_2_VITIS_LOOP_234_s_fu_180.fifo_conv_w_2_blk_n) begin
                            if (~AESL_inst_top.fifo_conv_w_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_conv_w_2_U' written by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_conv_w_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_conv_w_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_conv_w_2_U' read by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_conv_w_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertWeightToStream_U0.grp_ConvertWeightToStream_Pipeline_VITIS_LOOP_229_1_VITIS_LOOP_232_2_VITIS_LOOP_234_s_fu_180.fifo_conv_w_3_blk_n) begin
                            if (~AESL_inst_top.fifo_conv_w_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_conv_w_3_U' written by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_conv_w_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_conv_w_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_conv_w_3_U' read by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_conv_w_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertWeightToStream_U0.mode_c69_blk_n) begin
                            if (~AESL_inst_top.mode_c69_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.mode_c69_U' written by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c69_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.mode_c69_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.mode_c69_U' read by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c69_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    9: begin
                        if (~AESL_inst_top.ConvertWeightToStream_U0.grp_ConvertWeightToStream_Pipeline_VITIS_LOOP_251_5_VITIS_LOOP_254_6_VITIS_LOOP_257_s_fu_168.fifo_mm_w_blk_n) begin
                            if (~AESL_inst_top.fifo_mm_w_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_mm_w_U' written by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_mm_w_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_mm_w_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_mm_w_U' read by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_mm_w_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertWeightToStream_U0.mode_c68_blk_n) begin
                            if (~AESL_inst_top.mode_c68_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.mode_c68_U' written by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c68_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.mode_c68_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.mode_c68_U' read by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c68_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    0: begin
                        if (AESL_inst_top.ap_sync_ConvertWeightToStream_U0_ap_ready & AESL_inst_top.ConvertWeightToStream_U0.ap_idle & ~AESL_inst_top.ap_sync_entry_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'top.entry_proc_U0'");
                        end
                    end
                    1: begin
                        if (AESL_inst_top.ap_sync_ConvertWeightToStream_U0_ap_ready & AESL_inst_top.ConvertWeightToStream_U0.ap_idle & ~AESL_inst_top.ap_sync_Block_entry3_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'top.Block_entry3_proc_U0'");
                        end
                    end
                    2: begin
                        if (AESL_inst_top.ap_sync_ConvertWeightToStream_U0_ap_ready & AESL_inst_top.ConvertWeightToStream_U0.ap_idle & ~AESL_inst_top.ap_sync_ConvertBias_BN_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'top.ConvertBias_BN_U0'");
                        end
                    end
                    3: begin
                        if (AESL_inst_top.ap_sync_ConvertWeightToStream_U0_ap_ready & AESL_inst_top.ConvertWeightToStream_U0.ap_idle & ~AESL_inst_top.ap_sync_ConvertInputToStream_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'top.ConvertInputToStream_U0'");
                        end
                    end
                    endcase
                end
                8 : begin
                    case(index2)
                    7: begin
                        if (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.fifo_conv_w_blk_n) begin
                            if (~AESL_inst_top.fifo_conv_w_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_conv_w_U' written by process 'top.ConvertWeightToStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_conv_w_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_conv_w_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_conv_w_U' read by process 'top.ConvertWeightToStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_conv_w_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.fifo_conv_w_1_blk_n) begin
                            if (~AESL_inst_top.fifo_conv_w_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_conv_w_1_U' written by process 'top.ConvertWeightToStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_conv_w_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_conv_w_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_conv_w_1_U' read by process 'top.ConvertWeightToStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_conv_w_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.fifo_conv_w_2_blk_n) begin
                            if (~AESL_inst_top.fifo_conv_w_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_conv_w_2_U' written by process 'top.ConvertWeightToStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_conv_w_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_conv_w_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_conv_w_2_U' read by process 'top.ConvertWeightToStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_conv_w_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.fifo_conv_w_3_blk_n) begin
                            if (~AESL_inst_top.fifo_conv_w_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_conv_w_3_U' written by process 'top.ConvertWeightToStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_conv_w_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_conv_w_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_conv_w_3_U' read by process 'top.ConvertWeightToStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_conv_w_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvWeightToArray_U0.mode_blk_n) begin
                            if (~AESL_inst_top.mode_c69_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.mode_c69_U' written by process 'top.ConvertWeightToStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c69_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.mode_c69_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.mode_c69_U' read by process 'top.ConvertWeightToStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c69_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    10: begin
                        if (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.Conv_SA_W_blk_n) begin
                            if (~AESL_inst_top.Conv_SA_W_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Conv_SA_W_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Conv_SA_W_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Conv_SA_W_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.Conv_SA_W_1_blk_n) begin
                            if (~AESL_inst_top.Conv_SA_W_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Conv_SA_W_1_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Conv_SA_W_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Conv_SA_W_1_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.Conv_SA_W_2_blk_n) begin
                            if (~AESL_inst_top.Conv_SA_W_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Conv_SA_W_2_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Conv_SA_W_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Conv_SA_W_2_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.Conv_SA_W_3_blk_n) begin
                            if (~AESL_inst_top.Conv_SA_W_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Conv_SA_W_3_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Conv_SA_W_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Conv_SA_W_3_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.Conv_SA_W_4_blk_n) begin
                            if (~AESL_inst_top.Conv_SA_W_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Conv_SA_W_4_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Conv_SA_W_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Conv_SA_W_4_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.Conv_SA_W_5_blk_n) begin
                            if (~AESL_inst_top.Conv_SA_W_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Conv_SA_W_5_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Conv_SA_W_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Conv_SA_W_5_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.Conv_SA_W_6_blk_n) begin
                            if (~AESL_inst_top.Conv_SA_W_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Conv_SA_W_6_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Conv_SA_W_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Conv_SA_W_6_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.Conv_SA_W_7_blk_n) begin
                            if (~AESL_inst_top.Conv_SA_W_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Conv_SA_W_7_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Conv_SA_W_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Conv_SA_W_7_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.Conv_SA_W_8_blk_n) begin
                            if (~AESL_inst_top.Conv_SA_W_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Conv_SA_W_8_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Conv_SA_W_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Conv_SA_W_8_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.Conv_SA_W_9_blk_n) begin
                            if (~AESL_inst_top.Conv_SA_W_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Conv_SA_W_9_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Conv_SA_W_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Conv_SA_W_9_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.Conv_SA_W_10_blk_n) begin
                            if (~AESL_inst_top.Conv_SA_W_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Conv_SA_W_10_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Conv_SA_W_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Conv_SA_W_10_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.Conv_SA_W_11_blk_n) begin
                            if (~AESL_inst_top.Conv_SA_W_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Conv_SA_W_11_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Conv_SA_W_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Conv_SA_W_11_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.Conv_SA_W_12_blk_n) begin
                            if (~AESL_inst_top.Conv_SA_W_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Conv_SA_W_12_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Conv_SA_W_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Conv_SA_W_12_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.Conv_SA_W_13_blk_n) begin
                            if (~AESL_inst_top.Conv_SA_W_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Conv_SA_W_13_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Conv_SA_W_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Conv_SA_W_13_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.Conv_SA_W_14_blk_n) begin
                            if (~AESL_inst_top.Conv_SA_W_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Conv_SA_W_14_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Conv_SA_W_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Conv_SA_W_14_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvWeightToArray_U0.grp_ConvWeightToArray_Pipeline_VITIS_LOOP_275_1_VITIS_LOOP_278_2_fu_112.Conv_SA_W_15_blk_n) begin
                            if (~AESL_inst_top.Conv_SA_W_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Conv_SA_W_15_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Conv_SA_W_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Conv_SA_W_15_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvWeightToArray_U0.num_w_sa_loc_c_blk_n) begin
                            if (~AESL_inst_top.num_w_sa_loc_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.num_w_sa_loc_c_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.num_w_sa_loc_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.num_w_sa_loc_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.num_w_sa_loc_c_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.num_w_sa_loc_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvWeightToArray_U0.mode_c67_blk_n) begin
                            if (~AESL_inst_top.mode_c67_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.mode_c67_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c67_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.mode_c67_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.mode_c67_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c67_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.start_for_MuxWeightStream_U0_U.if_full_n & AESL_inst_top.ConvWeightToArray_U0.ap_start & ~AESL_inst_top.ConvWeightToArray_U0.real_start & (trans_in_cnt_1 == trans_out_cnt_1) & ~AESL_inst_top.start_for_MuxWeightStream_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'top.start_for_MuxWeightStream_U0_U' read by process 'top.MuxWeightStream_U0',");
                        end
                    end
                    1: begin
                        if (~AESL_inst_top.num_w_sa_loc_c36_channel_U.if_empty_n & AESL_inst_top.ConvWeightToArray_U0.ap_idle & ~AESL_inst_top.num_w_sa_loc_c36_channel_U.if_write) begin
                            if (~AESL_inst_top.num_w_sa_loc_c36_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.num_w_sa_loc_c36_channel_U' written by process 'top.Block_entry3_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.num_w_sa_loc_c36_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.num_w_sa_loc_c36_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.num_w_sa_loc_c36_channel_U' read by process 'top.Block_entry3_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.num_w_sa_loc_c36_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                9 : begin
                    case(index2)
                    7: begin
                        if (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.fifo_mm_w_blk_n) begin
                            if (~AESL_inst_top.fifo_mm_w_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_mm_w_U' written by process 'top.ConvertWeightToStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_mm_w_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_mm_w_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_mm_w_U' read by process 'top.ConvertWeightToStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_mm_w_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MMWeightToArray_U0.mode_blk_n) begin
                            if (~AESL_inst_top.mode_c68_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.mode_c68_U' written by process 'top.ConvertWeightToStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c68_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.mode_c68_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.mode_c68_U' read by process 'top.ConvertWeightToStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c68_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    10: begin
                        if (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.MM_SA_W_blk_n) begin
                            if (~AESL_inst_top.MM_SA_W_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_SA_W_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_SA_W_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_SA_W_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.MM_SA_W_1_blk_n) begin
                            if (~AESL_inst_top.MM_SA_W_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_SA_W_1_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_SA_W_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_SA_W_1_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.MM_SA_W_2_blk_n) begin
                            if (~AESL_inst_top.MM_SA_W_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_SA_W_2_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_SA_W_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_SA_W_2_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.MM_SA_W_3_blk_n) begin
                            if (~AESL_inst_top.MM_SA_W_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_SA_W_3_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_SA_W_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_SA_W_3_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.MM_SA_W_4_blk_n) begin
                            if (~AESL_inst_top.MM_SA_W_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_SA_W_4_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_SA_W_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_SA_W_4_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.MM_SA_W_5_blk_n) begin
                            if (~AESL_inst_top.MM_SA_W_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_SA_W_5_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_SA_W_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_SA_W_5_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.MM_SA_W_6_blk_n) begin
                            if (~AESL_inst_top.MM_SA_W_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_SA_W_6_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_SA_W_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_SA_W_6_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.MM_SA_W_7_blk_n) begin
                            if (~AESL_inst_top.MM_SA_W_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_SA_W_7_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_SA_W_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_SA_W_7_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.MM_SA_W_8_blk_n) begin
                            if (~AESL_inst_top.MM_SA_W_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_SA_W_8_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_SA_W_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_SA_W_8_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.MM_SA_W_9_blk_n) begin
                            if (~AESL_inst_top.MM_SA_W_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_SA_W_9_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_SA_W_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_SA_W_9_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.MM_SA_W_10_blk_n) begin
                            if (~AESL_inst_top.MM_SA_W_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_SA_W_10_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_SA_W_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_SA_W_10_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.MM_SA_W_11_blk_n) begin
                            if (~AESL_inst_top.MM_SA_W_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_SA_W_11_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_SA_W_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_SA_W_11_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.MM_SA_W_12_blk_n) begin
                            if (~AESL_inst_top.MM_SA_W_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_SA_W_12_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_SA_W_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_SA_W_12_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.MM_SA_W_13_blk_n) begin
                            if (~AESL_inst_top.MM_SA_W_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_SA_W_13_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_SA_W_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_SA_W_13_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.MM_SA_W_14_blk_n) begin
                            if (~AESL_inst_top.MM_SA_W_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_SA_W_14_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_SA_W_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_SA_W_14_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MMWeightToArray_U0.grp_MMWeightToArray_Pipeline_VITIS_LOOP_295_1_fu_78.MM_SA_W_15_blk_n) begin
                            if (~AESL_inst_top.MM_SA_W_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_SA_W_15_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_SA_W_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_SA_W_15_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    1: begin
                        if (~AESL_inst_top.num_w_sa_loc_c35_channel_U.if_empty_n & AESL_inst_top.MMWeightToArray_U0.ap_idle & ~AESL_inst_top.num_w_sa_loc_c35_channel_U.if_write) begin
                            if (~AESL_inst_top.num_w_sa_loc_c35_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.num_w_sa_loc_c35_channel_U' written by process 'top.Block_entry3_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.num_w_sa_loc_c35_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.num_w_sa_loc_c35_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.num_w_sa_loc_c35_channel_U' read by process 'top.Block_entry3_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.num_w_sa_loc_c35_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                10 : begin
                    case(index2)
                    8: begin
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.Conv_SA_W_blk_n) begin
                            if (~AESL_inst_top.Conv_SA_W_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Conv_SA_W_U' written by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Conv_SA_W_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Conv_SA_W_U' read by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.Conv_SA_W_1_blk_n) begin
                            if (~AESL_inst_top.Conv_SA_W_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Conv_SA_W_1_U' written by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Conv_SA_W_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Conv_SA_W_1_U' read by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.Conv_SA_W_2_blk_n) begin
                            if (~AESL_inst_top.Conv_SA_W_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Conv_SA_W_2_U' written by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Conv_SA_W_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Conv_SA_W_2_U' read by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.Conv_SA_W_3_blk_n) begin
                            if (~AESL_inst_top.Conv_SA_W_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Conv_SA_W_3_U' written by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Conv_SA_W_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Conv_SA_W_3_U' read by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.Conv_SA_W_4_blk_n) begin
                            if (~AESL_inst_top.Conv_SA_W_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Conv_SA_W_4_U' written by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Conv_SA_W_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Conv_SA_W_4_U' read by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.Conv_SA_W_5_blk_n) begin
                            if (~AESL_inst_top.Conv_SA_W_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Conv_SA_W_5_U' written by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Conv_SA_W_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Conv_SA_W_5_U' read by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.Conv_SA_W_6_blk_n) begin
                            if (~AESL_inst_top.Conv_SA_W_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Conv_SA_W_6_U' written by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Conv_SA_W_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Conv_SA_W_6_U' read by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.Conv_SA_W_7_blk_n) begin
                            if (~AESL_inst_top.Conv_SA_W_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Conv_SA_W_7_U' written by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Conv_SA_W_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Conv_SA_W_7_U' read by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.Conv_SA_W_8_blk_n) begin
                            if (~AESL_inst_top.Conv_SA_W_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Conv_SA_W_8_U' written by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Conv_SA_W_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Conv_SA_W_8_U' read by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.Conv_SA_W_9_blk_n) begin
                            if (~AESL_inst_top.Conv_SA_W_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Conv_SA_W_9_U' written by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Conv_SA_W_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Conv_SA_W_9_U' read by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.Conv_SA_W_10_blk_n) begin
                            if (~AESL_inst_top.Conv_SA_W_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Conv_SA_W_10_U' written by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Conv_SA_W_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Conv_SA_W_10_U' read by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.Conv_SA_W_11_blk_n) begin
                            if (~AESL_inst_top.Conv_SA_W_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Conv_SA_W_11_U' written by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Conv_SA_W_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Conv_SA_W_11_U' read by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.Conv_SA_W_12_blk_n) begin
                            if (~AESL_inst_top.Conv_SA_W_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Conv_SA_W_12_U' written by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Conv_SA_W_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Conv_SA_W_12_U' read by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.Conv_SA_W_13_blk_n) begin
                            if (~AESL_inst_top.Conv_SA_W_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Conv_SA_W_13_U' written by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Conv_SA_W_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Conv_SA_W_13_U' read by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.Conv_SA_W_14_blk_n) begin
                            if (~AESL_inst_top.Conv_SA_W_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Conv_SA_W_14_U' written by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Conv_SA_W_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Conv_SA_W_14_U' read by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.Conv_SA_W_15_blk_n) begin
                            if (~AESL_inst_top.Conv_SA_W_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Conv_SA_W_15_U' written by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Conv_SA_W_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Conv_SA_W_15_U' read by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Conv_SA_W_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.num_w_sa_loc_blk_n) begin
                            if (~AESL_inst_top.num_w_sa_loc_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.num_w_sa_loc_c_U' written by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.num_w_sa_loc_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.num_w_sa_loc_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.num_w_sa_loc_c_U' read by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.num_w_sa_loc_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.mode_blk_n) begin
                            if (~AESL_inst_top.mode_c67_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.mode_c67_U' written by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c67_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.mode_c67_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.mode_c67_U' read by process 'top.ConvWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c67_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.start_for_MuxWeightStream_U0_U.if_empty_n & AESL_inst_top.MuxWeightStream_U0.ap_idle & ~AESL_inst_top.start_for_MuxWeightStream_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'top.start_for_MuxWeightStream_U0_U' written by process 'top.ConvWeightToArray_U0',");
                        end
                    end
                    9: begin
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.MM_SA_W_blk_n) begin
                            if (~AESL_inst_top.MM_SA_W_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_SA_W_U' written by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_SA_W_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_SA_W_U' read by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.MM_SA_W_1_blk_n) begin
                            if (~AESL_inst_top.MM_SA_W_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_SA_W_1_U' written by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_SA_W_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_SA_W_1_U' read by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.MM_SA_W_2_blk_n) begin
                            if (~AESL_inst_top.MM_SA_W_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_SA_W_2_U' written by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_SA_W_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_SA_W_2_U' read by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.MM_SA_W_3_blk_n) begin
                            if (~AESL_inst_top.MM_SA_W_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_SA_W_3_U' written by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_SA_W_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_SA_W_3_U' read by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.MM_SA_W_4_blk_n) begin
                            if (~AESL_inst_top.MM_SA_W_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_SA_W_4_U' written by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_SA_W_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_SA_W_4_U' read by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.MM_SA_W_5_blk_n) begin
                            if (~AESL_inst_top.MM_SA_W_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_SA_W_5_U' written by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_SA_W_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_SA_W_5_U' read by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.MM_SA_W_6_blk_n) begin
                            if (~AESL_inst_top.MM_SA_W_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_SA_W_6_U' written by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_SA_W_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_SA_W_6_U' read by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.MM_SA_W_7_blk_n) begin
                            if (~AESL_inst_top.MM_SA_W_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_SA_W_7_U' written by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_SA_W_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_SA_W_7_U' read by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.MM_SA_W_8_blk_n) begin
                            if (~AESL_inst_top.MM_SA_W_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_SA_W_8_U' written by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_SA_W_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_SA_W_8_U' read by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.MM_SA_W_9_blk_n) begin
                            if (~AESL_inst_top.MM_SA_W_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_SA_W_9_U' written by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_SA_W_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_SA_W_9_U' read by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.MM_SA_W_10_blk_n) begin
                            if (~AESL_inst_top.MM_SA_W_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_SA_W_10_U' written by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_SA_W_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_SA_W_10_U' read by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.MM_SA_W_11_blk_n) begin
                            if (~AESL_inst_top.MM_SA_W_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_SA_W_11_U' written by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_SA_W_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_SA_W_11_U' read by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.MM_SA_W_12_blk_n) begin
                            if (~AESL_inst_top.MM_SA_W_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_SA_W_12_U' written by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_SA_W_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_SA_W_12_U' read by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.MM_SA_W_13_blk_n) begin
                            if (~AESL_inst_top.MM_SA_W_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_SA_W_13_U' written by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_SA_W_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_SA_W_13_U' read by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.MM_SA_W_14_blk_n) begin
                            if (~AESL_inst_top.MM_SA_W_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_SA_W_14_U' written by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_SA_W_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_SA_W_14_U' read by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.MM_SA_W_15_blk_n) begin
                            if (~AESL_inst_top.MM_SA_W_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_SA_W_15_U' written by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_SA_W_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_SA_W_15_U' read by process 'top.MMWeightToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_SA_W_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    11: begin
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.fifo_SA_W_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_W_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_W_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_W_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_W_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.fifo_SA_W_1_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_W_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_W_1_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_W_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_W_1_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.fifo_SA_W_2_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_W_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_W_2_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_W_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_W_2_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.fifo_SA_W_3_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_W_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_W_3_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_W_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_W_3_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.fifo_SA_W_4_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_W_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_W_4_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_W_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_W_4_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.fifo_SA_W_5_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_W_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_W_5_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_W_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_W_5_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.fifo_SA_W_6_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_W_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_W_6_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_W_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_W_6_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.fifo_SA_W_7_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_W_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_W_7_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_W_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_W_7_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.fifo_SA_W_8_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_W_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_W_8_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_W_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_W_8_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.fifo_SA_W_9_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_W_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_W_9_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_W_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_W_9_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.fifo_SA_W_10_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_W_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_W_10_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_W_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_W_10_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.fifo_SA_W_11_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_W_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_W_11_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_W_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_W_11_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.fifo_SA_W_12_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_W_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_W_12_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_W_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_W_12_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.fifo_SA_W_13_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_W_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_W_13_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_W_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_W_13_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.fifo_SA_W_14_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_W_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_W_14_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_W_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_W_14_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.MuxWeightStream_U0.grp_MuxWeightStream_Pipeline_VITIS_LOOP_314_1_fu_140.fifo_SA_W_15_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_W_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_W_15_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_W_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_W_15_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                11 : begin
                    case(index2)
                    6: begin
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_278.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_A_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_A_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_A_U' written by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_A_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_A_U' read by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_300.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_A_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_A_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_A_1_U' written by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_A_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_A_1_U' read by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_322.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_A_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_A_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_A_2_U' written by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_A_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_A_2_U' read by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_344.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_A_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_A_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_A_3_U' written by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_A_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_A_3_U' read by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_366.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_A_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_A_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_A_4_U' written by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_A_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_A_4_U' read by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_388.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_A_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_A_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_A_5_U' written by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_A_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_A_5_U' read by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_410.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_A_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_A_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_A_6_U' written by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_A_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_A_6_U' read by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_432.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_A_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_A_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_A_7_U' written by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_A_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_A_7_U' read by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_454.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_A_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_A_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_A_8_U' written by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_A_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_A_8_U' read by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_476.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_A_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_A_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_A_9_U' written by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_A_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_A_9_U' read by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_498.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_A_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_A_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_A_10_U' written by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_A_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_A_10_U' read by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_520.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_A_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_A_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_A_11_U' written by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_A_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_A_11_U' read by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_542.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_A_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_A_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_A_12_U' written by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_A_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_A_12_U' read by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_564.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_A_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_A_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_A_13_U' written by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_A_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_A_13_U' read by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_586.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_A_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_A_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_A_14_U' written by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_A_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_A_14_U' read by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_608.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_A_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_A_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_A_15_U' written by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_A_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_A_15_U' read by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_A_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.num_a_sa_2_loc_blk_n) begin
                            if (~AESL_inst_top.num_a_sa_2_loc_c42_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.num_a_sa_2_loc_c42_U' written by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.num_a_sa_2_loc_c42_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.num_a_sa_2_loc_c42_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.num_a_sa_2_loc_c42_U' read by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.num_a_sa_2_loc_c42_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.mode_blk_n) begin
                            if (~AESL_inst_top.mode_c66_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.mode_c66_U' written by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c66_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.mode_c66_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.mode_c66_U' read by process 'top.ConvertInputToArray_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c66_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    10: begin
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_278.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_W_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_W_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_W_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_W_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_W_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_300.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_W_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_W_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_W_1_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_W_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_W_1_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_322.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_W_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_W_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_W_2_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_W_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_W_2_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_344.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_W_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_W_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_W_3_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_W_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_W_3_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_366.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_W_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_W_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_W_4_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_W_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_W_4_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_388.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_W_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_W_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_W_5_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_W_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_W_5_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_410.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_W_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_W_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_W_6_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_W_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_W_6_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_432.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_W_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_W_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_W_7_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_W_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_W_7_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_454.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_W_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_W_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_W_8_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_W_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_W_8_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_476.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_W_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_W_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_W_9_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_W_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_W_9_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_498.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_W_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_W_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_W_10_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_W_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_W_10_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_520.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_W_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_W_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_W_11_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_W_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_W_11_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_542.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_W_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_W_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_W_12_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_W_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_W_12_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_564.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_W_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_W_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_W_13_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_W_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_W_13_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_586.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_W_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_W_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_W_14_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_W_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_W_14_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_608.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_W_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_W_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_W_15_U' written by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_W_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_W_15_U' read by process 'top.MuxWeightStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_W_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    12: begin
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_278.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_278.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_1_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_1_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_1_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_278.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_2_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_2_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_2_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_278.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_3_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_3_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_3_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_300.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_4_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_4_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_300.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_1_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_5_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_5_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_300.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_2_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_6_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_6_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_300.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_3_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_7_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_7_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_322.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_8_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_8_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_322.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_1_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_9_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_9_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_322.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_2_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_10_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_10_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_322.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_3_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_11_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_11_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_344.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_12_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_12_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_344.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_1_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_13_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_13_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_344.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_2_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_14_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_14_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_344.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_3_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_15_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_15_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_366.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_16_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_16_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_366.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_1_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_17_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_17_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_366.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_2_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_18_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_18_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_366.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_3_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_19_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_19_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_388.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_20_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_20_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_388.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_1_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_21_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_21_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_388.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_2_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_22_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_22_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_388.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_3_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_23_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_23_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_410.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_24_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_24_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_410.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_1_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_25_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_25_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_410.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_2_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_26_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_26_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_410.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_3_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_27_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_27_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_432.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_28_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_28_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_432.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_1_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_29_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_29_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_432.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_2_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_30_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_30_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_432.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_3_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_31_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_31_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_454.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_32_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_32_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_454.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_1_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_33_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_33_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_454.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_2_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_34_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_34_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_454.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_3_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_35_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_35_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_476.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_36_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_36_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_476.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_1_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_37_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_37_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_476.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_2_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_38_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_38_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_476.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_3_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_39_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_39_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_498.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_40_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_40_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_40_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_40_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_40_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_40_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_498.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_1_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_41_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_41_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_41_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_41_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_41_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_41_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_498.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_2_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_42_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_42_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_42_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_42_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_42_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_42_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_498.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_3_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_43_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_43_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_43_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_43_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_43_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_43_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_520.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_44_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_44_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_44_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_44_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_44_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_44_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_520.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_1_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_45_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_45_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_45_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_45_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_45_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_45_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_520.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_2_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_46_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_46_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_46_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_46_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_46_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_46_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_520.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_3_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_47_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_47_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_47_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_47_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_47_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_47_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_542.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_48_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_48_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_48_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_48_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_48_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_48_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_542.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_1_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_49_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_49_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_49_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_49_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_49_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_49_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_542.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_2_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_50_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_50_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_50_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_50_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_50_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_50_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_542.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_3_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_51_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_51_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_51_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_51_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_51_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_51_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_564.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_52_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_52_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_52_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_52_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_52_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_52_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_564.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_1_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_53_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_53_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_53_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_53_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_53_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_53_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_564.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_2_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_54_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_54_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_54_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_54_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_54_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_54_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_564.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_3_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_55_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_55_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_55_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_55_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_55_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_55_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_586.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_56_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_56_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_56_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_56_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_56_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_56_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_586.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_1_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_57_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_57_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_57_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_57_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_57_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_57_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_586.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_2_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_58_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_58_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_58_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_58_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_58_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_58_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_586.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_3_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_59_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_59_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_59_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_59_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_59_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_59_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_608.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_0_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_60_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_60_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_60_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_60_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_60_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_60_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_608.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_1_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_61_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_61_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_61_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_61_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_61_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_61_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_608.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_2_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_62_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_62_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_62_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_62_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_62_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_62_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.grp_PE_fu_608.grp_PE_Pipeline_VITIS_LOOP_385_5_fu_64.fifo_SA_O_0_0_3_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_63_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_63_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_63_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_63_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_63_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_63_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.num_a_sa_2_loc_c_blk_n) begin
                            if (~AESL_inst_top.num_a_sa_2_loc_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.num_a_sa_2_loc_c_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.num_a_sa_2_loc_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.num_a_sa_2_loc_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.num_a_sa_2_loc_c_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.num_a_sa_2_loc_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.Compute_U0.mode_c65_blk_n) begin
                            if (~AESL_inst_top.mode_c65_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.mode_c65_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c65_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.mode_c65_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.mode_c65_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c65_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    1: begin
                        if (~AESL_inst_top.out_c_1_loc_c41_channel_U.if_empty_n & AESL_inst_top.Compute_U0.ap_idle & ~AESL_inst_top.out_c_1_loc_c41_channel_U.if_write) begin
                            if (~AESL_inst_top.out_c_1_loc_c41_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.out_c_1_loc_c41_channel_U' written by process 'top.Block_entry3_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.out_c_1_loc_c41_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.out_c_1_loc_c41_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.out_c_1_loc_c41_channel_U' read by process 'top.Block_entry3_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.out_c_1_loc_c41_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    13: begin
                        if (~AESL_inst_top.Compute_U0.out_c_1_loc_c40_blk_n) begin
                            if (~AESL_inst_top.out_c_1_loc_c40_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.out_c_1_loc_c40_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.out_c_1_loc_c40_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.out_c_1_loc_c40_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.out_c_1_loc_c40_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.out_c_1_loc_c40_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                12 : begin
                    case(index2)
                    11: begin
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_1_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_1_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_1_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_2_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_2_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_2_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_3_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_3_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_3_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_4_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_4_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_4_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_5_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_5_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_5_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_6_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_6_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_6_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_7_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_7_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_7_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_8_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_8_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_8_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_9_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_9_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_9_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_10_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_10_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_10_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_11_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_11_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_11_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_12_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_12_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_12_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_13_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_13_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_13_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_14_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_14_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_14_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_15_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_15_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_15_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_16_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_16_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_16_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_17_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_17_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_17_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_18_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_18_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_18_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_19_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_19_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_19_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_20_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_20_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_20_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_21_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_21_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_21_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_22_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_22_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_22_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_23_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_23_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_23_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_24_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_24_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_24_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_25_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_25_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_25_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_26_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_26_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_26_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_27_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_27_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_27_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_28_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_28_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_28_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_29_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_29_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_29_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_30_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_30_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_30_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_31_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_31_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_31_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_32_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_32_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_32_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_33_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_33_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_33_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_34_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_34_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_34_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_35_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_35_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_35_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_36_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_36_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_36_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_37_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_37_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_37_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_38_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_38_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_38_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_39_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_39_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_39_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_40_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_40_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_40_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_40_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_40_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_40_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_40_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_41_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_41_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_41_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_41_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_41_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_41_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_41_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_42_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_42_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_42_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_42_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_42_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_42_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_42_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_43_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_43_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_43_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_43_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_43_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_43_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_43_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_44_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_44_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_44_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_44_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_44_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_44_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_44_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_45_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_45_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_45_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_45_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_45_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_45_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_45_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_46_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_46_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_46_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_46_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_46_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_46_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_46_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_47_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_47_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_47_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_47_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_47_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_47_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_47_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_48_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_48_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_48_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_48_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_48_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_48_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_48_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_49_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_49_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_49_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_49_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_49_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_49_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_49_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_50_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_50_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_50_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_50_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_50_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_50_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_50_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_51_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_51_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_51_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_51_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_51_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_51_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_51_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_52_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_52_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_52_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_52_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_52_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_52_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_52_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_53_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_53_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_53_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_53_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_53_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_53_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_53_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_54_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_54_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_54_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_54_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_54_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_54_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_54_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_55_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_55_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_55_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_55_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_55_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_55_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_55_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_56_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_56_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_56_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_56_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_56_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_56_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_56_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_57_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_57_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_57_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_57_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_57_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_57_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_57_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_58_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_58_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_58_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_58_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_58_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_58_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_58_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_59_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_59_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_59_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_59_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_59_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_59_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_59_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_60_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_60_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_60_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_60_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_60_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_60_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_60_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_61_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_61_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_61_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_61_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_61_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_61_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_61_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_62_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_62_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_62_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_62_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_62_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_62_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_62_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.fifo_SA_O_63_blk_n) begin
                            if (~AESL_inst_top.fifo_SA_O_63_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_SA_O_63_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_63_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_SA_O_63_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_SA_O_63_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_SA_O_63_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.num_a_sa_2_loc_blk_n) begin
                            if (~AESL_inst_top.num_a_sa_2_loc_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.num_a_sa_2_loc_c_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.num_a_sa_2_loc_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.num_a_sa_2_loc_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.num_a_sa_2_loc_c_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.num_a_sa_2_loc_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.mode_blk_n) begin
                            if (~AESL_inst_top.mode_c65_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.mode_c65_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c65_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.mode_c65_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.mode_c65_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c65_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    13: begin
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_570_1_fu_464.fifo_CONV3_ACC_blk_n) begin
                            if (~AESL_inst_top.fifo_CONV3_ACC_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_CONV3_ACC_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_CONV3_ACC_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_CONV3_ACC_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_570_1_fu_464.fifo_CONV3_ACC_1_blk_n) begin
                            if (~AESL_inst_top.fifo_CONV3_ACC_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_CONV3_ACC_1_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_CONV3_ACC_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_CONV3_ACC_1_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_570_1_fu_464.fifo_CONV3_ACC_2_blk_n) begin
                            if (~AESL_inst_top.fifo_CONV3_ACC_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_CONV3_ACC_2_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_CONV3_ACC_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_CONV3_ACC_2_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_570_1_fu_464.fifo_CONV3_ACC_3_blk_n) begin
                            if (~AESL_inst_top.fifo_CONV3_ACC_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_CONV3_ACC_3_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_CONV3_ACC_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_CONV3_ACC_3_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_570_1_fu_464.fifo_CONV3_ACC_4_blk_n) begin
                            if (~AESL_inst_top.fifo_CONV3_ACC_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_CONV3_ACC_4_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_CONV3_ACC_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_CONV3_ACC_4_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_570_1_fu_464.fifo_CONV3_ACC_5_blk_n) begin
                            if (~AESL_inst_top.fifo_CONV3_ACC_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_CONV3_ACC_5_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_CONV3_ACC_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_CONV3_ACC_5_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_570_1_fu_464.fifo_CONV3_ACC_6_blk_n) begin
                            if (~AESL_inst_top.fifo_CONV3_ACC_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_CONV3_ACC_6_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_CONV3_ACC_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_CONV3_ACC_6_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_570_1_fu_464.fifo_CONV3_ACC_7_blk_n) begin
                            if (~AESL_inst_top.fifo_CONV3_ACC_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_CONV3_ACC_7_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_CONV3_ACC_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_CONV3_ACC_7_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_570_1_fu_464.fifo_CONV3_ACC_8_blk_n) begin
                            if (~AESL_inst_top.fifo_CONV3_ACC_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_CONV3_ACC_8_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_CONV3_ACC_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_CONV3_ACC_8_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_570_1_fu_464.fifo_CONV3_ACC_9_blk_n) begin
                            if (~AESL_inst_top.fifo_CONV3_ACC_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_CONV3_ACC_9_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_CONV3_ACC_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_CONV3_ACC_9_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_570_1_fu_464.fifo_CONV3_ACC_10_blk_n) begin
                            if (~AESL_inst_top.fifo_CONV3_ACC_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_CONV3_ACC_10_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_CONV3_ACC_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_CONV3_ACC_10_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_570_1_fu_464.fifo_CONV3_ACC_11_blk_n) begin
                            if (~AESL_inst_top.fifo_CONV3_ACC_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_CONV3_ACC_11_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_CONV3_ACC_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_CONV3_ACC_11_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_570_1_fu_464.fifo_CONV3_ACC_12_blk_n) begin
                            if (~AESL_inst_top.fifo_CONV3_ACC_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_CONV3_ACC_12_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_CONV3_ACC_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_CONV3_ACC_12_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_570_1_fu_464.fifo_CONV3_ACC_13_blk_n) begin
                            if (~AESL_inst_top.fifo_CONV3_ACC_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_CONV3_ACC_13_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_CONV3_ACC_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_CONV3_ACC_13_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_570_1_fu_464.fifo_CONV3_ACC_14_blk_n) begin
                            if (~AESL_inst_top.fifo_CONV3_ACC_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_CONV3_ACC_14_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_CONV3_ACC_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_CONV3_ACC_14_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_570_1_fu_464.fifo_CONV3_ACC_15_blk_n) begin
                            if (~AESL_inst_top.fifo_CONV3_ACC_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_CONV3_ACC_15_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_CONV3_ACC_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_CONV3_ACC_15_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.N_c_blk_n) begin
                            if (~AESL_inst_top.N_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.N_c_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.N_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.N_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.N_c_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.N_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.mode_c64_blk_n) begin
                            if (~AESL_inst_top.mode_c64_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.mode_c64_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c64_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.mode_c64_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.mode_c64_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c64_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    16: begin
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.MM_OUT_blk_n) begin
                            if (~AESL_inst_top.MM_OUT_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_OUT_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_OUT_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_OUT_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.MM_OUT_1_blk_n) begin
                            if (~AESL_inst_top.MM_OUT_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_OUT_1_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_OUT_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_OUT_1_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.MM_OUT_2_blk_n) begin
                            if (~AESL_inst_top.MM_OUT_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_OUT_2_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_OUT_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_OUT_2_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.MM_OUT_3_blk_n) begin
                            if (~AESL_inst_top.MM_OUT_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_OUT_3_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_OUT_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_OUT_3_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.MM_OUT_4_blk_n) begin
                            if (~AESL_inst_top.MM_OUT_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_OUT_4_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_OUT_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_OUT_4_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.MM_OUT_5_blk_n) begin
                            if (~AESL_inst_top.MM_OUT_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_OUT_5_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_OUT_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_OUT_5_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.MM_OUT_6_blk_n) begin
                            if (~AESL_inst_top.MM_OUT_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_OUT_6_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_OUT_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_OUT_6_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.MM_OUT_7_blk_n) begin
                            if (~AESL_inst_top.MM_OUT_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_OUT_7_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_OUT_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_OUT_7_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.MM_OUT_8_blk_n) begin
                            if (~AESL_inst_top.MM_OUT_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_OUT_8_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_OUT_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_OUT_8_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.MM_OUT_9_blk_n) begin
                            if (~AESL_inst_top.MM_OUT_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_OUT_9_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_OUT_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_OUT_9_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.MM_OUT_10_blk_n) begin
                            if (~AESL_inst_top.MM_OUT_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_OUT_10_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_OUT_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_OUT_10_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.MM_OUT_11_blk_n) begin
                            if (~AESL_inst_top.MM_OUT_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_OUT_11_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_OUT_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_OUT_11_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.MM_OUT_12_blk_n) begin
                            if (~AESL_inst_top.MM_OUT_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_OUT_12_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_OUT_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_OUT_12_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.MM_OUT_13_blk_n) begin
                            if (~AESL_inst_top.MM_OUT_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_OUT_13_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_OUT_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_OUT_13_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.MM_OUT_14_blk_n) begin
                            if (~AESL_inst_top.MM_OUT_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_OUT_14_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_OUT_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_OUT_14_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.grp_ConvertToOutStream_Pipeline_VITIS_LOOP_592_5_VITIS_LOOP_595_6_VITIS_LOOP_598_7_V_fu_298.MM_OUT_15_blk_n) begin
                            if (~AESL_inst_top.MM_OUT_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_OUT_15_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_OUT_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_OUT_15_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.R_c_blk_n) begin
                            if (~AESL_inst_top.R_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.R_c_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.R_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.R_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.R_c_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.R_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    5: begin
                        if (~AESL_inst_top.ConvertToOutStream_U0.R_blk_n) begin
                            if (~AESL_inst_top.R_c44_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.R_c44_U' written by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.R_c44_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.R_c44_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.R_c44_U' read by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.R_c44_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvertToOutStream_U0.N_blk_n) begin
                            if (~AESL_inst_top.N_c49_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.N_c49_U' written by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.N_c49_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.N_c49_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.N_c49_U' read by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.N_c49_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.start_for_ConvertToOutStream_U0_U.if_empty_n & AESL_inst_top.ConvertToOutStream_U0.ap_idle & ~AESL_inst_top.start_for_ConvertToOutStream_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'top.start_for_ConvertToOutStream_U0_U' written by process 'top.Sliding_U0',");
                        end
                    end
                    endcase
                end
                13 : begin
                    case(index2)
                    12: begin
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.fifo_CONV3_ACC_blk_n) begin
                            if (~AESL_inst_top.fifo_CONV3_ACC_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_CONV3_ACC_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_CONV3_ACC_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_CONV3_ACC_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.fifo_CONV3_ACC_1_blk_n) begin
                            if (~AESL_inst_top.fifo_CONV3_ACC_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_CONV3_ACC_1_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_CONV3_ACC_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_CONV3_ACC_1_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.fifo_CONV3_ACC_2_blk_n) begin
                            if (~AESL_inst_top.fifo_CONV3_ACC_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_CONV3_ACC_2_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_CONV3_ACC_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_CONV3_ACC_2_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.fifo_CONV3_ACC_3_blk_n) begin
                            if (~AESL_inst_top.fifo_CONV3_ACC_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_CONV3_ACC_3_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_CONV3_ACC_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_CONV3_ACC_3_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.fifo_CONV3_ACC_4_blk_n) begin
                            if (~AESL_inst_top.fifo_CONV3_ACC_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_CONV3_ACC_4_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_CONV3_ACC_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_CONV3_ACC_4_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.fifo_CONV3_ACC_5_blk_n) begin
                            if (~AESL_inst_top.fifo_CONV3_ACC_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_CONV3_ACC_5_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_CONV3_ACC_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_CONV3_ACC_5_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.fifo_CONV3_ACC_6_blk_n) begin
                            if (~AESL_inst_top.fifo_CONV3_ACC_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_CONV3_ACC_6_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_CONV3_ACC_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_CONV3_ACC_6_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.fifo_CONV3_ACC_7_blk_n) begin
                            if (~AESL_inst_top.fifo_CONV3_ACC_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_CONV3_ACC_7_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_CONV3_ACC_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_CONV3_ACC_7_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.fifo_CONV3_ACC_8_blk_n) begin
                            if (~AESL_inst_top.fifo_CONV3_ACC_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_CONV3_ACC_8_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_CONV3_ACC_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_CONV3_ACC_8_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.fifo_CONV3_ACC_9_blk_n) begin
                            if (~AESL_inst_top.fifo_CONV3_ACC_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_CONV3_ACC_9_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_CONV3_ACC_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_CONV3_ACC_9_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.fifo_CONV3_ACC_10_blk_n) begin
                            if (~AESL_inst_top.fifo_CONV3_ACC_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_CONV3_ACC_10_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_CONV3_ACC_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_CONV3_ACC_10_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.fifo_CONV3_ACC_11_blk_n) begin
                            if (~AESL_inst_top.fifo_CONV3_ACC_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_CONV3_ACC_11_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_CONV3_ACC_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_CONV3_ACC_11_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.fifo_CONV3_ACC_12_blk_n) begin
                            if (~AESL_inst_top.fifo_CONV3_ACC_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_CONV3_ACC_12_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_CONV3_ACC_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_CONV3_ACC_12_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.fifo_CONV3_ACC_13_blk_n) begin
                            if (~AESL_inst_top.fifo_CONV3_ACC_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_CONV3_ACC_13_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_CONV3_ACC_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_CONV3_ACC_13_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.fifo_CONV3_ACC_14_blk_n) begin
                            if (~AESL_inst_top.fifo_CONV3_ACC_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_CONV3_ACC_14_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_CONV3_ACC_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_CONV3_ACC_14_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.fifo_CONV3_ACC_15_blk_n) begin
                            if (~AESL_inst_top.fifo_CONV3_ACC_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_CONV3_ACC_15_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_CONV3_ACC_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_CONV3_ACC_15_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_CONV3_ACC_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.N_blk_n) begin
                            if (~AESL_inst_top.N_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.N_c_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.N_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.N_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.N_c_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.N_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.mode_blk_n) begin
                            if (~AESL_inst_top.mode_c64_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.mode_c64_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c64_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.mode_c64_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.mode_c64_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c64_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    14: begin
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_1_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_1_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_1_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_2_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_2_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_2_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_3_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_3_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_3_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_4_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_4_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_4_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_5_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_5_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_5_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_6_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_6_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_6_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_7_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_7_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_7_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_8_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_8_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_8_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_9_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_9_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_9_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_10_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_10_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_10_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_11_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_11_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_11_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_12_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_12_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_12_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_13_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_13_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_13_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_14_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_14_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_14_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_15_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_15_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_15_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_16_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_16_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_16_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_17_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_17_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_17_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_18_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_18_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_18_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_19_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_19_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_19_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_20_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_20_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_20_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_21_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_21_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_21_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_22_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_22_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_22_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_23_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_23_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_23_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_24_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_24_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_24_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_25_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_25_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_25_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_26_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_26_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_26_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_27_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_27_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_27_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_28_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_28_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_28_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_29_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_29_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_29_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_30_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_30_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_30_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_31_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_31_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_31_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_32_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_32_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_32_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_33_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_33_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_33_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_34_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_34_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_34_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_35_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_35_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_35_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_36_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_36_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_36_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_37_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_37_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_37_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_38_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_38_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_38_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_39_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_39_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_39_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_40_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_40_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_40_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_40_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_40_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_40_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_40_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_41_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_41_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_41_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_41_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_41_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_41_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_41_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_42_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_42_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_42_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_42_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_42_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_42_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_42_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_43_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_43_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_43_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_43_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_43_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_43_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_43_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_44_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_44_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_44_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_44_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_44_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_44_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_44_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_45_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_45_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_45_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_45_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_45_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_45_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_45_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_46_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_46_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_46_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_46_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_46_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_46_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_46_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_47_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_47_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_47_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_47_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_47_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_47_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_47_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_48_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_48_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_48_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_48_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_48_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_48_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_48_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_49_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_49_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_49_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_49_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_49_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_49_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_49_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_50_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_50_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_50_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_50_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_50_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_50_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_50_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_51_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_51_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_51_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_51_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_51_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_51_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_51_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_52_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_52_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_52_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_52_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_52_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_52_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_52_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_53_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_53_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_53_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_53_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_53_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_53_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_53_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_54_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_54_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_54_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_54_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_54_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_54_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_54_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_55_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_55_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_55_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_55_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_55_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_55_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_55_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_56_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_56_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_56_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_56_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_56_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_56_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_56_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_57_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_57_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_57_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_57_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_57_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_57_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_57_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_58_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_58_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_58_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_58_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_58_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_58_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_58_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_59_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_59_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_59_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_59_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_59_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_59_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_59_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_60_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_60_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_60_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_60_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_60_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_60_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_60_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_61_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_61_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_61_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_61_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_61_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_61_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_61_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_62_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_62_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_62_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_62_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_62_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_62_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_62_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_63_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_63_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_63_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_63_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_63_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_63_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_63_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_64_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_64_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_64_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_64_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_64_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_64_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_64_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_65_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_65_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_65_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_65_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_65_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_65_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_65_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_66_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_66_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_66_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_66_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_66_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_66_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_66_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_67_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_67_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_67_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_67_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_67_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_67_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_67_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_68_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_68_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_68_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_68_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_68_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_68_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_68_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_69_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_69_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_69_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_69_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_69_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_69_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_69_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_70_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_70_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_70_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_70_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_70_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_70_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_70_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_71_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_71_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_71_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_71_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_71_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_71_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_71_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_72_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_72_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_72_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_72_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_72_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_72_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_72_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_73_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_73_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_73_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_73_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_73_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_73_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_73_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_74_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_74_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_74_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_74_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_74_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_74_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_74_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_75_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_75_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_75_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_75_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_75_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_75_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_75_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_76_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_76_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_76_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_76_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_76_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_76_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_76_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_77_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_77_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_77_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_77_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_77_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_77_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_77_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_78_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_78_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_78_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_78_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_78_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_78_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_78_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_79_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_79_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_79_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_79_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_79_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_79_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_79_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_80_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_80_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_80_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_80_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_80_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_80_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_80_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_81_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_81_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_81_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_81_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_81_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_81_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_81_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_82_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_82_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_82_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_82_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_82_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_82_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_82_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_83_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_83_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_83_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_83_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_83_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_83_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_83_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_84_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_84_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_84_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_84_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_84_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_84_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_84_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_85_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_85_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_85_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_85_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_85_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_85_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_85_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_86_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_86_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_86_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_86_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_86_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_86_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_86_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_87_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_87_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_87_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_87_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_87_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_87_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_87_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_88_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_88_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_88_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_88_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_88_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_88_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_88_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_89_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_89_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_89_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_89_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_89_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_89_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_89_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_90_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_90_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_90_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_90_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_90_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_90_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_90_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_91_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_91_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_91_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_91_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_91_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_91_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_91_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_92_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_92_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_92_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_92_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_92_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_92_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_92_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_93_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_93_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_93_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_93_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_93_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_93_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_93_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_94_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_94_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_94_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_94_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_94_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_94_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_94_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_95_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_95_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_95_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_95_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_95_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_95_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_95_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_96_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_96_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_96_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_96_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_96_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_96_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_96_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_97_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_97_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_97_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_97_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_97_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_97_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_97_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_98_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_98_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_98_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_98_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_98_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_98_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_98_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_99_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_99_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_99_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_99_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_99_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_99_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_99_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_100_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_100_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_100_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_100_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_100_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_100_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_100_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_101_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_101_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_101_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_101_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_101_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_101_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_101_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_102_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_102_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_102_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_102_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_102_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_102_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_102_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_103_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_103_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_103_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_103_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_103_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_103_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_103_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_104_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_104_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_104_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_104_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_104_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_104_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_104_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_105_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_105_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_105_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_105_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_105_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_105_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_105_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_106_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_106_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_106_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_106_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_106_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_106_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_106_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_107_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_107_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_107_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_107_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_107_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_107_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_107_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_108_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_108_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_108_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_108_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_108_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_108_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_108_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_109_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_109_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_109_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_109_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_109_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_109_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_109_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_110_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_110_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_110_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_110_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_110_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_110_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_110_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_111_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_111_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_111_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_111_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_111_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_111_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_111_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_112_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_112_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_112_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_112_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_112_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_112_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_112_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_113_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_113_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_113_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_113_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_113_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_113_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_113_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_114_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_114_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_114_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_114_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_114_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_114_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_114_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_115_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_115_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_115_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_115_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_115_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_115_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_115_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_116_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_116_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_116_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_116_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_116_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_116_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_116_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_117_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_117_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_117_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_117_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_117_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_117_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_117_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_118_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_118_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_118_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_118_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_118_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_118_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_118_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_119_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_119_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_119_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_119_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_119_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_119_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_119_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_120_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_120_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_120_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_120_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_120_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_120_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_120_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_121_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_121_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_121_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_121_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_121_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_121_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_121_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_122_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_122_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_122_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_122_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_122_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_122_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_122_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_123_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_123_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_123_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_123_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_123_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_123_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_123_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_124_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_124_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_124_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_124_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_124_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_124_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_124_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_125_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_125_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_125_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_125_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_125_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_125_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_125_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_126_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_126_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_126_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_126_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_126_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_126_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_126_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.grp_ConvToOutStream_Pipeline_VITIS_LOOP_624_1_VITIS_LOOP_627_2_VITIS_LOOP_630_3_VITI_fu_426.CONV3_OUT_127_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_127_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_127_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_127_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_127_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_127_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_127_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.out_r_1_loc_c37_blk_n) begin
                            if (~AESL_inst_top.out_r_1_loc_c37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.out_r_1_loc_c37_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.out_r_1_loc_c37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.out_r_1_loc_c37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.out_r_1_loc_c37_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.out_r_1_loc_c37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.out_c_1_loc_c39_blk_n) begin
                            if (~AESL_inst_top.out_c_1_loc_c39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.out_c_1_loc_c39_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.out_c_1_loc_c39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.out_c_1_loc_c39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.out_c_1_loc_c39_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.out_c_1_loc_c39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.M_c53_blk_n) begin
                            if (~AESL_inst_top.M_c53_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.M_c53_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.M_c53_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.M_c53_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.M_c53_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.M_c53_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.mode_c63_blk_n) begin
                            if (~AESL_inst_top.mode_c63_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.mode_c63_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c63_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.mode_c63_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.mode_c63_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c63_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    1: begin
                        if (~AESL_inst_top.out_r_1_loc_c38_channel_U.if_empty_n & AESL_inst_top.ConvToOutStream_U0.ap_idle & ~AESL_inst_top.out_r_1_loc_c38_channel_U.if_write) begin
                            if (~AESL_inst_top.out_r_1_loc_c38_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.out_r_1_loc_c38_channel_U' written by process 'top.Block_entry3_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.out_r_1_loc_c38_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.out_r_1_loc_c38_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.out_r_1_loc_c38_channel_U' read by process 'top.Block_entry3_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.out_r_1_loc_c38_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    11: begin
                        if (~AESL_inst_top.ConvToOutStream_U0.out_c_1_loc_blk_n) begin
                            if (~AESL_inst_top.out_c_1_loc_c40_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.out_c_1_loc_c40_U' written by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.out_c_1_loc_c40_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.out_c_1_loc_c40_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.out_c_1_loc_c40_U' read by process 'top.Compute_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.out_c_1_loc_c40_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    5: begin
                        if (~AESL_inst_top.ConvToOutStream_U0.M_blk_n) begin
                            if (~AESL_inst_top.M_c54_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.M_c54_U' written by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.M_c54_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.M_c54_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.M_c54_U' read by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.M_c54_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvToOutStream_U0.K_blk_n) begin
                            if (~AESL_inst_top.K_c57_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.K_c57_U' written by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.K_c57_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.K_c57_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.K_c57_U' read by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.K_c57_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    16: begin
                        if (~AESL_inst_top.ConvToOutStream_U0.K_c_blk_n) begin
                            if (~AESL_inst_top.K_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.K_c_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.K_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.K_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.K_c_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.K_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                14 : begin
                    case(index2)
                    13: begin
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_1_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_1_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_1_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_2_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_2_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_2_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_3_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_3_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_3_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_4_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_4_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_4_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_5_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_5_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_5_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_6_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_6_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_6_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_7_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_7_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_7_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_8_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_8_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_8_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_9_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_9_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_9_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_10_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_10_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_10_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_11_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_11_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_11_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_12_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_12_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_12_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_13_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_13_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_13_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_14_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_14_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_14_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_15_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_15_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_15_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_16_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_16_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_16_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_17_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_17_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_17_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_18_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_18_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_18_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_19_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_19_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_19_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_20_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_20_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_20_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_21_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_21_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_21_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_22_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_22_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_22_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_23_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_23_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_23_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_24_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_24_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_24_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_25_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_25_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_25_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_26_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_26_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_26_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_27_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_27_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_27_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_28_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_28_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_28_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_29_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_29_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_29_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_30_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_30_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_30_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_31_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_31_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_31_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_32_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_32_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_32_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_33_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_33_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_33_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_34_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_34_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_34_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_35_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_35_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_35_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_36_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_36_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_36_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_37_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_37_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_37_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_38_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_38_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_38_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_39_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_39_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_39_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_40_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_40_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_40_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_40_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_40_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_40_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_40_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_41_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_41_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_41_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_41_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_41_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_41_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_41_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_42_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_42_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_42_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_42_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_42_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_42_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_42_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_43_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_43_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_43_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_43_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_43_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_43_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_43_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_44_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_44_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_44_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_44_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_44_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_44_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_44_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_45_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_45_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_45_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_45_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_45_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_45_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_45_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_46_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_46_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_46_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_46_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_46_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_46_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_46_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_47_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_47_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_47_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_47_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_47_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_47_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_47_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_48_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_48_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_48_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_48_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_48_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_48_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_48_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_49_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_49_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_49_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_49_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_49_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_49_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_49_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_50_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_50_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_50_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_50_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_50_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_50_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_50_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_51_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_51_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_51_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_51_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_51_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_51_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_51_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_52_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_52_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_52_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_52_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_52_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_52_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_52_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_53_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_53_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_53_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_53_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_53_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_53_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_53_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_54_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_54_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_54_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_54_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_54_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_54_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_54_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_55_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_55_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_55_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_55_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_55_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_55_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_55_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_56_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_56_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_56_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_56_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_56_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_56_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_56_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_57_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_57_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_57_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_57_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_57_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_57_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_57_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_58_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_58_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_58_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_58_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_58_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_58_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_58_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_59_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_59_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_59_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_59_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_59_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_59_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_59_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_60_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_60_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_60_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_60_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_60_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_60_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_60_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_61_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_61_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_61_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_61_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_61_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_61_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_61_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_62_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_62_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_62_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_62_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_62_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_62_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_62_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_63_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_63_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_63_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_63_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_63_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_63_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_63_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_64_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_64_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_64_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_64_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_64_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_64_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_64_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_65_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_65_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_65_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_65_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_65_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_65_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_65_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_66_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_66_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_66_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_66_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_66_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_66_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_66_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_67_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_67_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_67_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_67_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_67_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_67_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_67_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_68_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_68_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_68_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_68_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_68_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_68_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_68_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_69_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_69_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_69_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_69_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_69_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_69_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_69_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_70_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_70_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_70_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_70_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_70_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_70_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_70_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_71_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_71_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_71_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_71_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_71_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_71_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_71_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_72_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_72_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_72_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_72_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_72_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_72_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_72_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_73_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_73_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_73_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_73_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_73_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_73_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_73_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_74_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_74_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_74_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_74_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_74_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_74_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_74_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_75_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_75_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_75_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_75_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_75_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_75_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_75_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_76_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_76_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_76_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_76_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_76_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_76_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_76_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_77_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_77_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_77_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_77_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_77_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_77_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_77_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_78_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_78_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_78_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_78_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_78_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_78_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_78_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_79_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_79_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_79_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_79_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_79_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_79_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_79_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_80_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_80_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_80_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_80_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_80_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_80_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_80_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_81_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_81_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_81_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_81_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_81_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_81_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_81_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_82_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_82_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_82_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_82_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_82_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_82_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_82_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_83_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_83_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_83_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_83_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_83_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_83_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_83_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_84_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_84_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_84_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_84_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_84_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_84_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_84_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_85_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_85_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_85_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_85_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_85_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_85_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_85_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_86_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_86_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_86_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_86_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_86_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_86_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_86_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_87_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_87_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_87_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_87_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_87_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_87_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_87_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_88_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_88_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_88_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_88_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_88_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_88_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_88_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_89_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_89_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_89_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_89_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_89_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_89_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_89_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_90_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_90_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_90_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_90_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_90_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_90_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_90_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_91_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_91_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_91_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_91_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_91_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_91_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_91_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_92_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_92_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_92_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_92_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_92_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_92_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_92_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_93_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_93_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_93_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_93_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_93_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_93_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_93_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_94_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_94_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_94_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_94_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_94_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_94_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_94_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_95_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_95_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_95_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_95_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_95_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_95_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_95_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_96_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_96_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_96_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_96_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_96_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_96_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_96_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_97_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_97_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_97_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_97_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_97_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_97_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_97_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_98_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_98_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_98_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_98_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_98_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_98_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_98_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_99_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_99_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_99_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_99_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_99_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_99_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_99_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_100_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_100_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_100_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_100_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_100_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_100_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_100_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_101_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_101_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_101_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_101_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_101_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_101_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_101_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_102_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_102_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_102_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_102_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_102_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_102_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_102_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_103_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_103_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_103_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_103_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_103_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_103_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_103_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_104_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_104_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_104_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_104_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_104_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_104_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_104_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_105_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_105_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_105_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_105_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_105_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_105_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_105_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_106_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_106_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_106_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_106_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_106_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_106_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_106_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_107_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_107_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_107_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_107_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_107_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_107_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_107_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_108_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_108_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_108_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_108_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_108_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_108_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_108_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_109_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_109_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_109_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_109_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_109_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_109_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_109_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_110_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_110_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_110_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_110_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_110_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_110_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_110_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_111_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_111_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_111_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_111_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_111_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_111_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_111_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_112_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_112_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_112_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_112_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_112_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_112_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_112_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_113_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_113_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_113_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_113_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_113_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_113_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_113_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_114_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_114_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_114_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_114_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_114_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_114_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_114_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_115_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_115_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_115_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_115_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_115_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_115_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_115_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_116_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_116_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_116_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_116_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_116_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_116_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_116_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_117_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_117_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_117_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_117_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_117_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_117_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_117_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_118_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_118_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_118_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_118_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_118_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_118_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_118_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_119_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_119_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_119_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_119_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_119_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_119_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_119_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_120_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_120_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_120_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_120_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_120_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_120_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_120_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_121_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_121_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_121_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_121_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_121_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_121_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_121_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_122_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_122_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_122_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_122_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_122_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_122_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_122_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_123_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_123_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_123_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_123_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_123_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_123_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_123_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_124_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_124_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_124_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_124_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_124_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_124_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_124_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_125_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_125_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_125_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_125_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_125_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_125_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_125_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_126_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_126_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_126_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_126_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_126_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_126_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_126_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_OUT_127_blk_n) begin
                            if (~AESL_inst_top.CONV3_OUT_127_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_OUT_127_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_127_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_OUT_127_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_OUT_127_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_OUT_127_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.out_r_1_loc_blk_n) begin
                            if (~AESL_inst_top.out_r_1_loc_c37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.out_r_1_loc_c37_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.out_r_1_loc_c37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.out_r_1_loc_c37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.out_r_1_loc_c37_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.out_r_1_loc_c37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.out_c_1_loc_blk_n) begin
                            if (~AESL_inst_top.out_c_1_loc_c39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.out_c_1_loc_c39_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.out_c_1_loc_c39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.out_c_1_loc_c39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.out_c_1_loc_c39_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.out_c_1_loc_c39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.M_blk_n) begin
                            if (~AESL_inst_top.M_c53_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.M_c53_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.M_c53_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.M_c53_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.M_c53_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.M_c53_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.mode_blk_n) begin
                            if (~AESL_inst_top.mode_c63_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.mode_c63_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c63_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.mode_c63_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.mode_c63_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c63_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    2: begin
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_1_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_1_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_1_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_2_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_2_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_2_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_3_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_3_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_3_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_4_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_4_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_4_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_5_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_5_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_5_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_6_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_6_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_6_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_7_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_7_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_7_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_8_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_8_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_8_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_9_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_9_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_9_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_10_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_10_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_10_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_11_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_11_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_11_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_12_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_12_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_12_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_13_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_13_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_13_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_14_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_14_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_14_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_15_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_15_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_15_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_16_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_16_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_16_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_17_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_17_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_17_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_18_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_18_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_18_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_19_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_19_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_19_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_20_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_20_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_20_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_21_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_21_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_21_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_22_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_22_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_22_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_23_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_23_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_23_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_24_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_24_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_24_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_25_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_25_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_25_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_26_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_26_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_26_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_27_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_27_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_27_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_28_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_28_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_28_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_29_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_29_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_29_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_30_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_30_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_30_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_31_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_31_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_31_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_32_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_32_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_32_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_33_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_33_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_33_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_34_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_34_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_34_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_35_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_35_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_35_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_36_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_36_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_36_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_37_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_37_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_37_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_38_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_38_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_38_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_39_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_39_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_39_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_40_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_40_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_40_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_40_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_40_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_40_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_40_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_41_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_41_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_41_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_41_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_41_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_41_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_41_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_42_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_42_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_42_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_42_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_42_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_42_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_42_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_43_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_43_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_43_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_43_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_43_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_43_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_43_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_44_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_44_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_44_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_44_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_44_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_44_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_44_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_45_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_45_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_45_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_45_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_45_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_45_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_45_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_46_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_46_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_46_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_46_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_46_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_46_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_46_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_47_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_47_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_47_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_47_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_47_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_47_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_47_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_48_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_48_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_48_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_48_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_48_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_48_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_48_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_49_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_49_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_49_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_49_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_49_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_49_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_49_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_50_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_50_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_50_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_50_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_50_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_50_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_50_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_51_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_51_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_51_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_51_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_51_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_51_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_51_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_52_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_52_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_52_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_52_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_52_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_52_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_52_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_53_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_53_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_53_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_53_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_53_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_53_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_53_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_54_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_54_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_54_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_54_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_54_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_54_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_54_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_55_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_55_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_55_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_55_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_55_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_55_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_55_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_56_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_56_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_56_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_56_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_56_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_56_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_56_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_57_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_57_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_57_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_57_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_57_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_57_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_57_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_58_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_58_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_58_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_58_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_58_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_58_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_58_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_59_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_59_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_59_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_59_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_59_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_59_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_59_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_60_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_60_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_60_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_60_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_60_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_60_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_60_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_61_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_61_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_61_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_61_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_61_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_61_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_61_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_62_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_62_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_62_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_62_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_62_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_62_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_62_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_63_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_63_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_63_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_63_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_63_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_63_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_63_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_64_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_64_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_64_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_64_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_64_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_64_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_64_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_65_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_65_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_65_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_65_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_65_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_65_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_65_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_66_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_66_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_66_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_66_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_66_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_66_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_66_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_67_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_67_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_67_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_67_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_67_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_67_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_67_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_68_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_68_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_68_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_68_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_68_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_68_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_68_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_69_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_69_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_69_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_69_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_69_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_69_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_69_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_70_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_70_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_70_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_70_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_70_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_70_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_70_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_71_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_71_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_71_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_71_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_71_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_71_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_71_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_72_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_72_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_72_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_72_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_72_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_72_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_72_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_73_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_73_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_73_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_73_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_73_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_73_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_73_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_74_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_74_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_74_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_74_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_74_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_74_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_74_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_75_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_75_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_75_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_75_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_75_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_75_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_75_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_76_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_76_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_76_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_76_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_76_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_76_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_76_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_77_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_77_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_77_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_77_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_77_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_77_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_77_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_78_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_78_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_78_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_78_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_78_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_78_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_78_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_79_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_79_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_79_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_79_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_79_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_79_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_79_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_80_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_80_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_80_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_80_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_80_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_80_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_80_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_81_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_81_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_81_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_81_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_81_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_81_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_81_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_82_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_82_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_82_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_82_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_82_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_82_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_82_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_83_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_83_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_83_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_83_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_83_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_83_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_83_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_84_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_84_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_84_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_84_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_84_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_84_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_84_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_85_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_85_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_85_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_85_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_85_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_85_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_85_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_86_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_86_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_86_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_86_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_86_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_86_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_86_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_87_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_87_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_87_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_87_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_87_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_87_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_87_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_88_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_88_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_88_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_88_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_88_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_88_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_88_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_89_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_89_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_89_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_89_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_89_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_89_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_89_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_90_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_90_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_90_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_90_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_90_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_90_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_90_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_91_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_91_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_91_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_91_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_91_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_91_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_91_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_92_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_92_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_92_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_92_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_92_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_92_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_92_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_93_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_93_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_93_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_93_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_93_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_93_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_93_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_94_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_94_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_94_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_94_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_94_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_94_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_94_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_95_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_95_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_95_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_95_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_95_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_95_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_95_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_96_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_96_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_96_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_96_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_96_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_96_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_96_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_97_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_97_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_97_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_97_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_97_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_97_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_97_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_98_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_98_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_98_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_98_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_98_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_98_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_98_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_99_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_99_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_99_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_99_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_99_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_99_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_99_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_100_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_100_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_100_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_100_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_100_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_100_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_100_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_101_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_101_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_101_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_101_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_101_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_101_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_101_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_102_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_102_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_102_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_102_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_102_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_102_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_102_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_103_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_103_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_103_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_103_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_103_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_103_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_103_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_104_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_104_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_104_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_104_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_104_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_104_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_104_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_105_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_105_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_105_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_105_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_105_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_105_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_105_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_106_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_106_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_106_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_106_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_106_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_106_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_106_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_107_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_107_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_107_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_107_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_107_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_107_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_107_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_108_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_108_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_108_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_108_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_108_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_108_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_108_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_109_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_109_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_109_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_109_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_109_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_109_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_109_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_110_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_110_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_110_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_110_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_110_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_110_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_110_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_111_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_111_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_111_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_111_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_111_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_111_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_111_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_112_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_112_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_112_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_112_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_112_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_112_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_112_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_113_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_113_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_113_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_113_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_113_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_113_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_113_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_114_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_114_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_114_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_114_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_114_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_114_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_114_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_115_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_115_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_115_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_115_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_115_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_115_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_115_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_116_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_116_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_116_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_116_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_116_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_116_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_116_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_117_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_117_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_117_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_117_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_117_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_117_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_117_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_118_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_118_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_118_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_118_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_118_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_118_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_118_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_119_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_119_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_119_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_119_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_119_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_119_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_119_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_120_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_120_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_120_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_120_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_120_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_120_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_120_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_121_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_121_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_121_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_121_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_121_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_121_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_121_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_122_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_122_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_122_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_122_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_122_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_122_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_122_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_123_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_123_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_123_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_123_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_123_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_123_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_123_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_124_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_124_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_124_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_124_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_124_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_124_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_124_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_125_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_125_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_125_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_125_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_125_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_125_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_125_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_126_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_126_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_126_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_126_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_126_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_126_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_126_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.fifo_bias_127_blk_n) begin
                            if (~AESL_inst_top.fifo_bias_127_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_bias_127_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_127_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_bias_127_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_bias_127_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_bias_127_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.start_for_ConvBias_U0_U.if_empty_n & AESL_inst_top.ConvBias_U0.ap_idle & ~AESL_inst_top.start_for_ConvBias_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'top.start_for_ConvBias_U0_U' written by process 'top.ConvertBias_BN_U0',");
                        end
                    end
                    15: begin
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_1_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_1_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_1_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_2_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_2_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_2_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_3_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_3_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_3_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_4_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_4_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_4_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_5_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_5_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_5_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_6_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_6_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_6_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_7_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_7_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_7_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_8_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_8_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_8_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_9_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_9_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_9_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_10_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_10_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_10_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_11_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_11_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_11_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_12_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_12_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_12_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_13_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_13_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_13_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_14_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_14_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_14_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_15_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_15_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_15_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_16_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_16_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_16_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_17_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_17_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_17_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_18_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_18_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_18_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_19_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_19_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_19_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_20_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_20_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_20_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_21_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_21_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_21_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_22_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_22_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_22_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_23_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_23_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_23_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_24_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_24_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_24_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_25_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_25_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_25_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_26_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_26_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_26_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_27_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_27_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_27_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_28_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_28_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_28_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_29_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_29_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_29_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_30_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_30_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_30_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_31_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_31_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_31_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_32_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_32_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_32_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_33_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_33_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_33_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_34_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_34_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_34_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_35_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_35_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_35_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_36_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_36_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_36_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_37_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_37_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_37_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_38_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_38_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_38_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_39_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_39_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_39_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_40_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_40_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_40_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_40_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_40_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_40_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_40_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_41_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_41_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_41_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_41_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_41_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_41_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_41_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_42_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_42_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_42_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_42_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_42_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_42_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_42_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_43_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_43_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_43_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_43_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_43_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_43_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_43_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_44_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_44_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_44_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_44_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_44_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_44_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_44_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_45_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_45_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_45_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_45_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_45_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_45_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_45_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_46_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_46_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_46_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_46_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_46_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_46_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_46_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_47_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_47_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_47_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_47_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_47_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_47_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_47_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_48_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_48_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_48_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_48_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_48_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_48_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_48_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_49_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_49_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_49_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_49_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_49_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_49_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_49_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_50_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_50_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_50_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_50_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_50_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_50_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_50_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_51_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_51_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_51_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_51_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_51_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_51_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_51_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_52_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_52_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_52_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_52_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_52_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_52_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_52_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_53_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_53_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_53_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_53_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_53_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_53_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_53_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_54_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_54_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_54_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_54_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_54_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_54_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_54_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_55_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_55_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_55_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_55_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_55_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_55_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_55_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_56_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_56_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_56_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_56_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_56_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_56_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_56_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_57_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_57_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_57_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_57_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_57_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_57_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_57_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_58_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_58_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_58_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_58_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_58_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_58_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_58_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_59_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_59_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_59_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_59_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_59_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_59_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_59_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_60_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_60_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_60_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_60_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_60_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_60_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_60_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_61_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_61_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_61_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_61_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_61_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_61_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_61_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_62_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_62_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_62_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_62_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_62_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_62_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_62_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_63_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_63_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_63_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_63_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_63_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_63_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_63_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_64_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_64_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_64_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_64_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_64_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_64_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_64_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_65_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_65_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_65_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_65_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_65_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_65_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_65_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_66_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_66_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_66_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_66_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_66_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_66_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_66_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_67_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_67_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_67_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_67_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_67_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_67_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_67_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_68_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_68_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_68_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_68_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_68_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_68_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_68_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_69_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_69_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_69_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_69_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_69_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_69_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_69_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_70_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_70_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_70_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_70_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_70_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_70_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_70_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_71_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_71_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_71_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_71_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_71_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_71_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_71_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_72_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_72_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_72_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_72_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_72_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_72_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_72_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_73_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_73_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_73_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_73_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_73_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_73_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_73_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_74_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_74_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_74_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_74_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_74_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_74_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_74_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_75_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_75_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_75_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_75_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_75_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_75_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_75_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_76_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_76_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_76_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_76_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_76_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_76_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_76_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_77_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_77_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_77_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_77_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_77_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_77_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_77_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_78_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_78_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_78_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_78_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_78_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_78_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_78_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_79_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_79_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_79_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_79_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_79_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_79_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_79_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_80_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_80_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_80_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_80_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_80_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_80_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_80_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_81_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_81_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_81_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_81_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_81_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_81_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_81_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_82_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_82_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_82_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_82_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_82_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_82_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_82_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_83_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_83_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_83_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_83_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_83_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_83_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_83_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_84_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_84_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_84_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_84_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_84_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_84_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_84_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_85_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_85_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_85_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_85_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_85_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_85_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_85_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_86_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_86_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_86_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_86_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_86_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_86_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_86_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_87_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_87_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_87_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_87_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_87_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_87_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_87_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_88_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_88_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_88_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_88_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_88_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_88_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_88_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_89_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_89_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_89_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_89_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_89_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_89_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_89_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_90_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_90_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_90_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_90_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_90_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_90_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_90_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_91_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_91_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_91_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_91_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_91_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_91_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_91_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_92_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_92_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_92_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_92_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_92_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_92_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_92_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_93_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_93_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_93_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_93_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_93_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_93_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_93_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_94_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_94_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_94_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_94_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_94_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_94_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_94_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_95_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_95_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_95_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_95_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_95_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_95_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_95_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_96_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_96_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_96_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_96_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_96_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_96_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_96_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_97_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_97_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_97_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_97_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_97_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_97_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_97_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_98_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_98_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_98_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_98_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_98_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_98_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_98_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_99_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_99_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_99_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_99_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_99_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_99_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_99_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_100_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_100_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_100_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_100_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_100_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_100_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_100_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_101_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_101_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_101_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_101_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_101_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_101_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_101_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_102_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_102_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_102_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_102_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_102_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_102_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_102_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_103_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_103_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_103_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_103_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_103_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_103_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_103_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_104_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_104_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_104_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_104_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_104_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_104_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_104_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_105_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_105_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_105_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_105_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_105_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_105_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_105_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_106_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_106_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_106_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_106_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_106_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_106_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_106_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_107_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_107_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_107_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_107_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_107_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_107_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_107_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_108_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_108_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_108_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_108_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_108_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_108_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_108_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_109_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_109_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_109_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_109_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_109_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_109_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_109_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_110_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_110_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_110_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_110_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_110_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_110_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_110_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_111_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_111_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_111_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_111_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_111_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_111_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_111_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_112_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_112_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_112_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_112_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_112_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_112_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_112_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_113_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_113_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_113_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_113_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_113_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_113_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_113_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_114_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_114_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_114_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_114_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_114_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_114_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_114_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_115_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_115_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_115_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_115_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_115_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_115_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_115_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_116_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_116_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_116_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_116_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_116_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_116_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_116_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_117_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_117_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_117_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_117_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_117_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_117_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_117_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_118_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_118_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_118_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_118_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_118_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_118_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_118_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_119_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_119_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_119_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_119_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_119_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_119_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_119_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_120_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_120_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_120_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_120_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_120_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_120_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_120_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_121_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_121_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_121_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_121_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_121_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_121_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_121_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_122_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_122_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_122_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_122_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_122_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_122_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_122_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_123_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_123_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_123_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_123_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_123_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_123_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_123_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_124_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_124_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_124_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_124_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_124_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_124_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_124_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_125_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_125_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_125_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_125_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_125_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_125_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_125_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_126_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_126_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_126_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_126_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_126_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_126_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_126_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.grp_ConvBias_Pipeline_VITIS_LOOP_663_1_VITIS_LOOP_666_2_VITIS_LOOP_668_3_VITIS_LOOP_s_fu_886.CONV3_BIAS_127_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_127_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_127_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_127_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_127_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_127_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_127_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.out_r_1_loc_c_blk_n) begin
                            if (~AESL_inst_top.out_r_1_loc_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.out_r_1_loc_c_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.out_r_1_loc_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.out_r_1_loc_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.out_r_1_loc_c_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.out_r_1_loc_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.out_c_1_loc_c_blk_n) begin
                            if (~AESL_inst_top.out_c_1_loc_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.out_c_1_loc_c_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.out_c_1_loc_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.out_c_1_loc_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.out_c_1_loc_c_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.out_c_1_loc_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.M_c52_blk_n) begin
                            if (~AESL_inst_top.M_c52_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.M_c52_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.M_c52_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.M_c52_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.M_c52_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.M_c52_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBias_U0.mode_c62_blk_n) begin
                            if (~AESL_inst_top.mode_c62_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.mode_c62_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c62_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.mode_c62_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.mode_c62_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c62_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                15 : begin
                    case(index2)
                    14: begin
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_1_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_1_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_1_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_2_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_2_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_2_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_3_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_3_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_3_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_4_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_4_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_4_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_5_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_5_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_5_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_6_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_6_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_6_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_7_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_7_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_7_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_8_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_8_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_8_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_9_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_9_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_9_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_10_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_10_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_10_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_11_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_11_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_11_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_12_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_12_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_12_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_13_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_13_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_13_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_14_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_14_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_14_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_15_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_15_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_15_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_16_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_16_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_16_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_17_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_17_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_17_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_18_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_18_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_18_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_19_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_19_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_19_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_20_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_20_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_20_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_21_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_21_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_21_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_22_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_22_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_22_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_23_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_23_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_23_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_24_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_24_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_24_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_25_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_25_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_25_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_26_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_26_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_26_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_27_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_27_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_27_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_28_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_28_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_28_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_29_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_29_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_29_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_30_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_30_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_30_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_31_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_31_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_31_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_32_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_32_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_32_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_33_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_33_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_33_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_34_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_34_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_34_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_35_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_35_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_35_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_36_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_36_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_36_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_37_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_37_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_37_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_38_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_38_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_38_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_39_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_39_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_39_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_40_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_40_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_40_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_40_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_40_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_40_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_40_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_41_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_41_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_41_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_41_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_41_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_41_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_41_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_42_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_42_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_42_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_42_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_42_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_42_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_42_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_43_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_43_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_43_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_43_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_43_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_43_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_43_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_44_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_44_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_44_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_44_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_44_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_44_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_44_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_45_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_45_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_45_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_45_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_45_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_45_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_45_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_46_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_46_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_46_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_46_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_46_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_46_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_46_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_47_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_47_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_47_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_47_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_47_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_47_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_47_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_48_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_48_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_48_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_48_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_48_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_48_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_48_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_49_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_49_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_49_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_49_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_49_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_49_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_49_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_50_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_50_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_50_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_50_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_50_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_50_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_50_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_51_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_51_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_51_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_51_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_51_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_51_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_51_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_52_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_52_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_52_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_52_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_52_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_52_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_52_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_53_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_53_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_53_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_53_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_53_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_53_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_53_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_54_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_54_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_54_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_54_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_54_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_54_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_54_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_55_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_55_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_55_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_55_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_55_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_55_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_55_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_56_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_56_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_56_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_56_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_56_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_56_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_56_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_57_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_57_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_57_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_57_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_57_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_57_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_57_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_58_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_58_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_58_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_58_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_58_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_58_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_58_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_59_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_59_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_59_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_59_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_59_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_59_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_59_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_60_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_60_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_60_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_60_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_60_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_60_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_60_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_61_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_61_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_61_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_61_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_61_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_61_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_61_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_62_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_62_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_62_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_62_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_62_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_62_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_62_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_63_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_63_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_63_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_63_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_63_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_63_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_63_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_64_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_64_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_64_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_64_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_64_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_64_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_64_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_65_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_65_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_65_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_65_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_65_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_65_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_65_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_66_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_66_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_66_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_66_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_66_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_66_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_66_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_67_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_67_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_67_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_67_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_67_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_67_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_67_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_68_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_68_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_68_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_68_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_68_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_68_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_68_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_69_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_69_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_69_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_69_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_69_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_69_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_69_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_70_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_70_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_70_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_70_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_70_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_70_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_70_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_71_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_71_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_71_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_71_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_71_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_71_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_71_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_72_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_72_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_72_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_72_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_72_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_72_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_72_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_73_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_73_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_73_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_73_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_73_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_73_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_73_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_74_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_74_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_74_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_74_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_74_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_74_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_74_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_75_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_75_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_75_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_75_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_75_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_75_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_75_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_76_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_76_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_76_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_76_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_76_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_76_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_76_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_77_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_77_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_77_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_77_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_77_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_77_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_77_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_78_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_78_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_78_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_78_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_78_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_78_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_78_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_79_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_79_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_79_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_79_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_79_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_79_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_79_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_80_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_80_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_80_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_80_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_80_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_80_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_80_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_81_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_81_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_81_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_81_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_81_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_81_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_81_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_82_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_82_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_82_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_82_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_82_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_82_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_82_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_83_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_83_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_83_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_83_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_83_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_83_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_83_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_84_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_84_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_84_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_84_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_84_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_84_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_84_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_85_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_85_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_85_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_85_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_85_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_85_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_85_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_86_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_86_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_86_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_86_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_86_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_86_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_86_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_87_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_87_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_87_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_87_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_87_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_87_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_87_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_88_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_88_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_88_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_88_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_88_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_88_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_88_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_89_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_89_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_89_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_89_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_89_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_89_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_89_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_90_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_90_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_90_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_90_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_90_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_90_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_90_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_91_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_91_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_91_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_91_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_91_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_91_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_91_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_92_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_92_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_92_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_92_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_92_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_92_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_92_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_93_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_93_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_93_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_93_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_93_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_93_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_93_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_94_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_94_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_94_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_94_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_94_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_94_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_94_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_95_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_95_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_95_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_95_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_95_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_95_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_95_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_96_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_96_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_96_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_96_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_96_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_96_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_96_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_97_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_97_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_97_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_97_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_97_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_97_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_97_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_98_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_98_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_98_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_98_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_98_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_98_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_98_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_99_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_99_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_99_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_99_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_99_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_99_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_99_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_100_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_100_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_100_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_100_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_100_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_100_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_100_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_101_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_101_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_101_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_101_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_101_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_101_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_101_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_102_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_102_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_102_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_102_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_102_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_102_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_102_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_103_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_103_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_103_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_103_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_103_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_103_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_103_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_104_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_104_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_104_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_104_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_104_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_104_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_104_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_105_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_105_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_105_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_105_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_105_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_105_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_105_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_106_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_106_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_106_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_106_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_106_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_106_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_106_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_107_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_107_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_107_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_107_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_107_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_107_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_107_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_108_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_108_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_108_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_108_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_108_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_108_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_108_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_109_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_109_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_109_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_109_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_109_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_109_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_109_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_110_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_110_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_110_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_110_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_110_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_110_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_110_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_111_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_111_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_111_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_111_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_111_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_111_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_111_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_112_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_112_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_112_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_112_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_112_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_112_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_112_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_113_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_113_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_113_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_113_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_113_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_113_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_113_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_114_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_114_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_114_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_114_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_114_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_114_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_114_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_115_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_115_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_115_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_115_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_115_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_115_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_115_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_116_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_116_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_116_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_116_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_116_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_116_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_116_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_117_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_117_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_117_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_117_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_117_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_117_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_117_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_118_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_118_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_118_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_118_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_118_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_118_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_118_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_119_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_119_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_119_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_119_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_119_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_119_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_119_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_120_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_120_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_120_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_120_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_120_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_120_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_120_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_121_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_121_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_121_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_121_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_121_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_121_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_121_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_122_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_122_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_122_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_122_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_122_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_122_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_122_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_123_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_123_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_123_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_123_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_123_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_123_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_123_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_124_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_124_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_124_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_124_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_124_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_124_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_124_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_125_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_125_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_125_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_125_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_125_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_125_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_125_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_126_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_126_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_126_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_126_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_126_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_126_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_126_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_BIAS_127_blk_n) begin
                            if (~AESL_inst_top.CONV3_BIAS_127_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_BIAS_127_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_127_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_BIAS_127_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_BIAS_127_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_BIAS_127_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.out_r_1_loc_blk_n) begin
                            if (~AESL_inst_top.out_r_1_loc_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.out_r_1_loc_c_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.out_r_1_loc_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.out_r_1_loc_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.out_r_1_loc_c_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.out_r_1_loc_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.out_c_1_loc_blk_n) begin
                            if (~AESL_inst_top.out_c_1_loc_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.out_c_1_loc_c_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.out_c_1_loc_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.out_c_1_loc_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.out_c_1_loc_c_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.out_c_1_loc_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.M_blk_n) begin
                            if (~AESL_inst_top.M_c52_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.M_c52_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.M_c52_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.M_c52_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.M_c52_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.M_c52_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.mode_blk_n) begin
                            if (~AESL_inst_top.mode_c62_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.mode_c62_U' written by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c62_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.mode_c62_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.mode_c62_U' read by process 'top.ConvBias_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c62_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    16: begin
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_1_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_1_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_1_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_2_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_2_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_2_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_3_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_3_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_3_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_4_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_4_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_4_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_5_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_5_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_5_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_6_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_6_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_6_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_7_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_7_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_7_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_8_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_8_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_8_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_9_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_9_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_9_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_10_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_10_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_10_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_11_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_11_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_11_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_12_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_12_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_12_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_13_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_13_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_13_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_14_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_14_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_14_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_15_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_15_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_15_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_16_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_16_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_16_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_17_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_17_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_17_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_18_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_18_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_18_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_19_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_19_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_19_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_20_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_20_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_20_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_21_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_21_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_21_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_22_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_22_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_22_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_23_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_23_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_23_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_24_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_24_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_24_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_25_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_25_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_25_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_26_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_26_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_26_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_27_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_27_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_27_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_28_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_28_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_28_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_29_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_29_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_29_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_30_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_30_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_30_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_31_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_31_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_31_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_32_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_32_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_32_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_33_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_33_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_33_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_34_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_34_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_34_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_35_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_35_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_35_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_36_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_36_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_36_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_37_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_37_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_37_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_38_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_38_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_38_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_39_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_39_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_39_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_40_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_40_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_40_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_40_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_40_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_40_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_40_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_41_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_41_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_41_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_41_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_41_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_41_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_41_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_42_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_42_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_42_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_42_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_42_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_42_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_42_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_43_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_43_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_43_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_43_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_43_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_43_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_43_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_44_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_44_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_44_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_44_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_44_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_44_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_44_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_45_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_45_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_45_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_45_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_45_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_45_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_45_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_46_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_46_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_46_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_46_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_46_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_46_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_46_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_47_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_47_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_47_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_47_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_47_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_47_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_47_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_48_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_48_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_48_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_48_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_48_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_48_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_48_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_49_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_49_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_49_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_49_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_49_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_49_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_49_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_50_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_50_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_50_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_50_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_50_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_50_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_50_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_51_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_51_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_51_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_51_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_51_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_51_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_51_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_52_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_52_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_52_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_52_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_52_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_52_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_52_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_53_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_53_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_53_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_53_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_53_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_53_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_53_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_54_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_54_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_54_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_54_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_54_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_54_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_54_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_55_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_55_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_55_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_55_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_55_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_55_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_55_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_56_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_56_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_56_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_56_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_56_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_56_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_56_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_57_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_57_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_57_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_57_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_57_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_57_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_57_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_58_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_58_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_58_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_58_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_58_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_58_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_58_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_59_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_59_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_59_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_59_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_59_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_59_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_59_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_60_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_60_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_60_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_60_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_60_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_60_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_60_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_61_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_61_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_61_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_61_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_61_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_61_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_61_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_62_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_62_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_62_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_62_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_62_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_62_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_62_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_63_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_63_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_63_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_63_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_63_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_63_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_63_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_64_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_64_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_64_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_64_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_64_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_64_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_64_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_65_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_65_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_65_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_65_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_65_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_65_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_65_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_66_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_66_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_66_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_66_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_66_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_66_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_66_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_67_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_67_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_67_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_67_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_67_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_67_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_67_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_68_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_68_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_68_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_68_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_68_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_68_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_68_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_69_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_69_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_69_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_69_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_69_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_69_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_69_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_70_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_70_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_70_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_70_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_70_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_70_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_70_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_71_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_71_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_71_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_71_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_71_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_71_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_71_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_72_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_72_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_72_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_72_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_72_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_72_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_72_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_73_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_73_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_73_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_73_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_73_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_73_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_73_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_74_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_74_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_74_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_74_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_74_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_74_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_74_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_75_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_75_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_75_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_75_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_75_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_75_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_75_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_76_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_76_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_76_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_76_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_76_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_76_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_76_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_77_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_77_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_77_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_77_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_77_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_77_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_77_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_78_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_78_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_78_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_78_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_78_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_78_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_78_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_79_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_79_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_79_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_79_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_79_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_79_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_79_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_80_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_80_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_80_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_80_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_80_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_80_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_80_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_81_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_81_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_81_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_81_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_81_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_81_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_81_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_82_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_82_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_82_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_82_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_82_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_82_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_82_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_83_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_83_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_83_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_83_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_83_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_83_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_83_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_84_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_84_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_84_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_84_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_84_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_84_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_84_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_85_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_85_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_85_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_85_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_85_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_85_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_85_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_86_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_86_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_86_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_86_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_86_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_86_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_86_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_87_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_87_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_87_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_87_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_87_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_87_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_87_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_88_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_88_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_88_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_88_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_88_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_88_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_88_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_89_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_89_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_89_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_89_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_89_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_89_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_89_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_90_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_90_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_90_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_90_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_90_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_90_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_90_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_91_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_91_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_91_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_91_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_91_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_91_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_91_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_92_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_92_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_92_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_92_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_92_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_92_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_92_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_93_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_93_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_93_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_93_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_93_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_93_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_93_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_94_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_94_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_94_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_94_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_94_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_94_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_94_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_95_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_95_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_95_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_95_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_95_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_95_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_95_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_96_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_96_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_96_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_96_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_96_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_96_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_96_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_97_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_97_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_97_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_97_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_97_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_97_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_97_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_98_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_98_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_98_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_98_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_98_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_98_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_98_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_99_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_99_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_99_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_99_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_99_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_99_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_99_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_100_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_100_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_100_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_100_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_100_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_100_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_100_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_101_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_101_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_101_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_101_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_101_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_101_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_101_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_102_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_102_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_102_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_102_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_102_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_102_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_102_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_103_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_103_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_103_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_103_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_103_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_103_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_103_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_104_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_104_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_104_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_104_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_104_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_104_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_104_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_105_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_105_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_105_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_105_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_105_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_105_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_105_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_106_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_106_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_106_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_106_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_106_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_106_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_106_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_107_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_107_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_107_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_107_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_107_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_107_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_107_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_108_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_108_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_108_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_108_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_108_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_108_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_108_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_109_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_109_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_109_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_109_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_109_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_109_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_109_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_110_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_110_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_110_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_110_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_110_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_110_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_110_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_111_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_111_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_111_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_111_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_111_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_111_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_111_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_112_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_112_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_112_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_112_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_112_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_112_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_112_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_113_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_113_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_113_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_113_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_113_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_113_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_113_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_114_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_114_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_114_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_114_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_114_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_114_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_114_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_115_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_115_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_115_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_115_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_115_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_115_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_115_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_116_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_116_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_116_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_116_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_116_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_116_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_116_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_117_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_117_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_117_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_117_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_117_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_117_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_117_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_118_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_118_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_118_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_118_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_118_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_118_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_118_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_119_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_119_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_119_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_119_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_119_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_119_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_119_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_120_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_120_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_120_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_120_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_120_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_120_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_120_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_121_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_121_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_121_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_121_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_121_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_121_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_121_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_122_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_122_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_122_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_122_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_122_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_122_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_122_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_123_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_123_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_123_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_123_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_123_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_123_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_123_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_124_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_124_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_124_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_124_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_124_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_124_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_124_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_125_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_125_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_125_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_125_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_125_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_125_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_125_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_126_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_126_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_126_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_126_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_126_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_126_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_126_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.CONV3_NORM_127_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_127_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_127_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_127_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_127_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_127_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_127_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.M_c_blk_n) begin
                            if (~AESL_inst_top.M_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.M_c_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.M_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.M_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.M_c_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.M_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.mode_c_blk_n) begin
                            if (~AESL_inst_top.mode_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.mode_c_U' written by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.mode_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.mode_c_U' read by process 'top.ResOutput_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    2: begin
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_1_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_1_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_1_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_2_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_2_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_2_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_3_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_3_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_3_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_4_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_4_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_4_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_5_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_5_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_5_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_6_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_6_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_6_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_7_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_7_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_7_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_8_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_8_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_8_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_9_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_9_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_9_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_10_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_10_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_10_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_11_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_11_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_11_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_12_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_12_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_12_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_13_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_13_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_13_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_14_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_14_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_14_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_15_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_15_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_15_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_16_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_16_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_16_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_17_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_17_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_17_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_18_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_18_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_18_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_19_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_19_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_19_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_20_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_20_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_20_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_21_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_21_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_21_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_22_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_22_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_22_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_23_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_23_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_23_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_24_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_24_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_24_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_25_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_25_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_25_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_26_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_26_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_26_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_27_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_27_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_27_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_28_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_28_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_28_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_29_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_29_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_29_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_30_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_30_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_30_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_31_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_31_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_31_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_32_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_32_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_32_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_33_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_33_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_33_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_34_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_34_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_34_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_35_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_35_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_35_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_36_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_36_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_36_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_37_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_37_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_37_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_38_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_38_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_38_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_39_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_39_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_39_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_40_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_40_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_40_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_40_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_40_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_40_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_40_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_41_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_41_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_41_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_41_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_41_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_41_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_41_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_42_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_42_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_42_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_42_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_42_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_42_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_42_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_43_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_43_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_43_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_43_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_43_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_43_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_43_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_44_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_44_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_44_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_44_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_44_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_44_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_44_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_45_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_45_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_45_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_45_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_45_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_45_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_45_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_46_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_46_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_46_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_46_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_46_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_46_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_46_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_47_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_47_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_47_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_47_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_47_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_47_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_47_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_48_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_48_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_48_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_48_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_48_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_48_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_48_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_49_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_49_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_49_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_49_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_49_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_49_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_49_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_50_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_50_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_50_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_50_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_50_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_50_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_50_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_51_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_51_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_51_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_51_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_51_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_51_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_51_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_52_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_52_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_52_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_52_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_52_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_52_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_52_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_53_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_53_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_53_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_53_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_53_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_53_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_53_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_54_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_54_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_54_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_54_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_54_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_54_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_54_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_55_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_55_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_55_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_55_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_55_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_55_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_55_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_56_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_56_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_56_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_56_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_56_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_56_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_56_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_57_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_57_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_57_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_57_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_57_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_57_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_57_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_58_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_58_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_58_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_58_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_58_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_58_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_58_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_59_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_59_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_59_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_59_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_59_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_59_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_59_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_60_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_60_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_60_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_60_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_60_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_60_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_60_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_61_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_61_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_61_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_61_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_61_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_61_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_61_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_62_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_62_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_62_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_62_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_62_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_62_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_62_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_63_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_63_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_63_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_63_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_63_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_63_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_63_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_64_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_64_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_64_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_64_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_64_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_64_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_64_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_65_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_65_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_65_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_65_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_65_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_65_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_65_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_66_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_66_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_66_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_66_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_66_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_66_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_66_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_67_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_67_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_67_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_67_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_67_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_67_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_67_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_68_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_68_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_68_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_68_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_68_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_68_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_68_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_69_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_69_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_69_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_69_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_69_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_69_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_69_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_70_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_70_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_70_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_70_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_70_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_70_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_70_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_71_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_71_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_71_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_71_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_71_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_71_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_71_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_72_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_72_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_72_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_72_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_72_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_72_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_72_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_73_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_73_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_73_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_73_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_73_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_73_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_73_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_74_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_74_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_74_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_74_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_74_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_74_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_74_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_75_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_75_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_75_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_75_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_75_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_75_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_75_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_76_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_76_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_76_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_76_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_76_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_76_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_76_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_77_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_77_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_77_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_77_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_77_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_77_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_77_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_78_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_78_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_78_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_78_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_78_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_78_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_78_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_79_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_79_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_79_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_79_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_79_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_79_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_79_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_80_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_80_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_80_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_80_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_80_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_80_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_80_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_81_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_81_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_81_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_81_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_81_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_81_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_81_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_82_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_82_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_82_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_82_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_82_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_82_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_82_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_83_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_83_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_83_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_83_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_83_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_83_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_83_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_84_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_84_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_84_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_84_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_84_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_84_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_84_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_85_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_85_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_85_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_85_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_85_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_85_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_85_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_86_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_86_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_86_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_86_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_86_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_86_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_86_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_87_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_87_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_87_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_87_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_87_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_87_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_87_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_88_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_88_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_88_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_88_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_88_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_88_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_88_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_89_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_89_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_89_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_89_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_89_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_89_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_89_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_90_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_90_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_90_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_90_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_90_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_90_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_90_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_91_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_91_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_91_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_91_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_91_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_91_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_91_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_92_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_92_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_92_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_92_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_92_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_92_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_92_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_93_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_93_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_93_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_93_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_93_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_93_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_93_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_94_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_94_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_94_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_94_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_94_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_94_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_94_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_95_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_95_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_95_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_95_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_95_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_95_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_95_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_96_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_96_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_96_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_96_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_96_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_96_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_96_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_97_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_97_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_97_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_97_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_97_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_97_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_97_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_98_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_98_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_98_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_98_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_98_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_98_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_98_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_99_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_99_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_99_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_99_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_99_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_99_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_99_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_100_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_100_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_100_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_100_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_100_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_100_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_100_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_101_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_101_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_101_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_101_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_101_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_101_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_101_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_102_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_102_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_102_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_102_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_102_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_102_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_102_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_103_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_103_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_103_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_103_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_103_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_103_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_103_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_104_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_104_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_104_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_104_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_104_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_104_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_104_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_105_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_105_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_105_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_105_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_105_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_105_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_105_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_106_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_106_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_106_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_106_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_106_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_106_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_106_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_107_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_107_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_107_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_107_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_107_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_107_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_107_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_108_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_108_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_108_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_108_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_108_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_108_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_108_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_109_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_109_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_109_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_109_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_109_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_109_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_109_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_110_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_110_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_110_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_110_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_110_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_110_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_110_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_111_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_111_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_111_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_111_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_111_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_111_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_111_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_112_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_112_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_112_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_112_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_112_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_112_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_112_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_113_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_113_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_113_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_113_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_113_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_113_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_113_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_114_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_114_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_114_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_114_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_114_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_114_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_114_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_115_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_115_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_115_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_115_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_115_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_115_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_115_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_116_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_116_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_116_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_116_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_116_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_116_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_116_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_117_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_117_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_117_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_117_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_117_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_117_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_117_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_118_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_118_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_118_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_118_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_118_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_118_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_118_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_119_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_119_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_119_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_119_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_119_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_119_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_119_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_120_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_120_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_120_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_120_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_120_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_120_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_120_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_121_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_121_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_121_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_121_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_121_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_121_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_121_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_122_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_122_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_122_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_122_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_122_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_122_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_122_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_123_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_123_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_123_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_123_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_123_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_123_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_123_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_124_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_124_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_124_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_124_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_124_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_124_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_124_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_125_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_125_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_125_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_125_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_125_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_125_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_125_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_126_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_126_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_126_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_126_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_126_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_126_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_126_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ConvBN_U0.grp_ConvBN_Pipeline_VITIS_LOOP_688_1_VITIS_LOOP_691_2_fu_852.fifo_norm_127_blk_n) begin
                            if (~AESL_inst_top.fifo_norm_127_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.fifo_norm_127_U' written by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_127_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.fifo_norm_127_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.fifo_norm_127_U' read by process 'top.ConvertBias_BN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.fifo_norm_127_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.start_for_ConvBN_U0_U.if_empty_n & AESL_inst_top.ConvBN_U0.ap_idle & ~AESL_inst_top.start_for_ConvBN_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'top.start_for_ConvBN_U0_U' written by process 'top.ConvertBias_BN_U0',");
                        end
                    end
                    endcase
                end
                16 : begin
                    case(index2)
                    15: begin
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_0_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_1_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_1_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_1_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_2_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_2_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_2_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_3_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_3_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_3_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_4_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_4_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_4_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_5_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_5_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_5_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_6_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_6_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_6_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_7_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_7_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_7_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_8_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_8_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_8_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_9_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_9_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_9_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_10_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_10_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_10_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_11_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_11_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_11_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_12_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_12_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_12_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_13_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_13_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_13_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_14_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_14_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_14_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_15_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_15_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_15_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_16_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_16_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_16_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_17_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_17_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_17_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_18_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_18_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_18_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_19_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_19_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_19_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_20_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_20_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_20_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_21_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_21_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_21_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_22_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_22_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_22_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_23_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_23_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_23_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_24_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_24_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_24_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_25_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_25_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_25_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_26_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_26_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_26_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_27_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_27_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_27_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_28_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_28_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_28_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_29_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_29_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_29_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_30_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_30_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_30_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_31_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_31_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_31_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_32_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_32_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_32_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_33_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_33_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_33_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_34_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_34_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_34_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_35_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_35_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_35_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_36_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_36_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_36_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_37_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_37_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_37_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_38_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_38_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_38_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_39_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_39_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_39_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_40_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_40_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_40_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_40_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_40_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_40_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_40_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_41_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_41_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_41_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_41_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_41_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_41_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_41_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_42_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_42_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_42_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_42_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_42_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_42_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_42_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_43_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_43_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_43_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_43_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_43_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_43_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_43_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_44_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_44_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_44_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_44_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_44_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_44_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_44_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_45_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_45_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_45_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_45_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_45_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_45_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_45_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_46_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_46_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_46_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_46_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_46_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_46_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_46_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_47_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_47_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_47_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_47_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_47_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_47_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_47_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_48_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_48_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_48_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_48_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_48_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_48_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_48_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_49_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_49_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_49_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_49_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_49_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_49_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_49_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_50_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_50_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_50_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_50_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_50_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_50_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_50_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_51_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_51_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_51_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_51_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_51_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_51_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_51_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_52_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_52_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_52_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_52_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_52_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_52_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_52_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_53_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_53_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_53_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_53_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_53_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_53_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_53_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_54_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_54_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_54_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_54_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_54_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_54_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_54_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_55_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_55_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_55_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_55_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_55_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_55_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_55_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_56_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_56_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_56_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_56_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_56_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_56_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_56_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_57_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_57_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_57_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_57_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_57_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_57_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_57_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_58_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_58_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_58_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_58_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_58_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_58_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_58_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_59_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_59_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_59_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_59_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_59_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_59_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_59_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_60_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_60_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_60_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_60_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_60_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_60_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_60_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_61_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_61_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_61_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_61_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_61_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_61_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_61_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_62_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_62_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_62_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_62_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_62_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_62_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_62_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_63_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_63_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_63_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_63_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_63_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_63_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_63_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_64_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_64_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_64_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_64_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_64_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_64_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_64_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_65_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_65_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_65_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_65_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_65_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_65_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_65_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_66_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_66_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_66_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_66_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_66_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_66_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_66_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_67_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_67_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_67_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_67_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_67_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_67_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_67_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_68_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_68_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_68_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_68_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_68_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_68_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_68_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_69_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_69_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_69_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_69_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_69_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_69_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_69_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_70_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_70_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_70_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_70_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_70_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_70_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_70_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_71_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_71_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_71_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_71_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_71_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_71_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_71_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_72_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_72_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_72_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_72_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_72_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_72_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_72_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_73_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_73_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_73_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_73_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_73_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_73_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_73_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_74_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_74_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_74_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_74_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_74_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_74_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_74_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_75_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_75_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_75_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_75_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_75_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_75_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_75_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_76_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_76_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_76_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_76_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_76_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_76_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_76_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_77_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_77_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_77_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_77_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_77_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_77_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_77_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_78_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_78_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_78_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_78_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_78_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_78_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_78_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_79_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_79_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_79_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_79_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_79_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_79_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_79_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_80_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_80_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_80_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_80_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_80_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_80_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_80_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_81_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_81_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_81_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_81_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_81_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_81_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_81_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_82_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_82_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_82_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_82_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_82_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_82_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_82_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_83_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_83_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_83_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_83_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_83_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_83_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_83_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_84_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_84_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_84_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_84_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_84_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_84_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_84_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_85_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_85_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_85_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_85_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_85_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_85_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_85_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_86_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_86_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_86_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_86_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_86_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_86_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_86_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_87_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_87_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_87_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_87_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_87_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_87_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_87_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_88_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_88_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_88_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_88_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_88_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_88_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_88_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_89_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_89_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_89_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_89_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_89_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_89_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_89_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_90_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_90_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_90_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_90_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_90_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_90_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_90_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_91_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_91_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_91_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_91_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_91_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_91_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_91_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_92_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_92_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_92_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_92_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_92_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_92_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_92_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_93_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_93_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_93_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_93_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_93_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_93_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_93_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_94_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_94_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_94_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_94_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_94_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_94_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_94_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_95_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_95_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_95_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_95_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_95_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_95_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_95_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_96_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_96_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_96_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_96_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_96_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_96_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_96_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_97_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_97_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_97_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_97_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_97_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_97_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_97_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_98_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_98_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_98_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_98_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_98_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_98_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_98_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_99_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_99_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_99_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_99_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_99_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_99_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_99_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_100_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_100_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_100_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_100_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_100_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_100_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_100_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_101_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_101_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_101_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_101_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_101_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_101_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_101_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_102_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_102_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_102_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_102_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_102_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_102_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_102_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_103_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_103_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_103_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_103_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_103_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_103_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_103_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_104_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_104_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_104_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_104_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_104_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_104_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_104_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_105_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_105_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_105_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_105_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_105_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_105_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_105_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_106_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_106_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_106_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_106_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_106_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_106_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_106_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_107_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_107_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_107_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_107_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_107_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_107_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_107_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_108_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_108_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_108_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_108_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_108_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_108_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_108_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_109_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_109_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_109_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_109_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_109_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_109_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_109_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_110_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_110_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_110_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_110_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_110_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_110_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_110_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_111_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_111_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_111_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_111_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_111_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_111_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_111_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_112_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_112_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_112_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_112_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_112_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_112_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_112_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_113_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_113_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_113_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_113_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_113_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_113_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_113_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_114_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_114_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_114_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_114_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_114_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_114_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_114_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_115_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_115_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_115_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_115_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_115_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_115_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_115_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_116_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_116_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_116_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_116_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_116_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_116_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_116_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_117_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_117_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_117_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_117_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_117_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_117_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_117_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_118_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_118_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_118_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_118_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_118_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_118_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_118_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_119_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_119_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_119_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_119_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_119_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_119_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_119_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_120_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_120_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_120_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_120_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_120_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_120_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_120_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_121_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_121_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_121_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_121_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_121_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_121_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_121_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_122_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_122_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_122_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_122_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_122_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_122_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_122_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_123_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_123_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_123_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_123_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_123_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_123_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_123_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_124_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_124_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_124_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_124_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_124_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_124_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_124_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_125_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_125_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_125_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_125_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_125_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_125_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_125_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_126_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_126_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_126_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_126_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_126_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_126_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_126_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_718_1_VITIS_LOOP_721_2_VITIS_LOOP_724_3_fu_448.CONV3_NORM_127_blk_n) begin
                            if (~AESL_inst_top.CONV3_NORM_127_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.CONV3_NORM_127_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_127_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.CONV3_NORM_127_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.CONV3_NORM_127_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.CONV3_NORM_127_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.M_blk_n) begin
                            if (~AESL_inst_top.M_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.M_c_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.M_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.M_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.M_c_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.M_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.mode_blk_n) begin
                            if (~AESL_inst_top.mode_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.mode_c_U' written by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.mode_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.mode_c_U' read by process 'top.ConvBN_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.mode_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    12: begin
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_734_4_VITIS_LOOP_737_5_VITIS_LOOP_740_6_VITIS_LOOP_fu_406.MM_OUT_0_blk_n) begin
                            if (~AESL_inst_top.MM_OUT_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_OUT_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_OUT_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_OUT_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_734_4_VITIS_LOOP_737_5_VITIS_LOOP_740_6_VITIS_LOOP_fu_406.MM_OUT_1_blk_n) begin
                            if (~AESL_inst_top.MM_OUT_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_OUT_1_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_OUT_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_OUT_1_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_734_4_VITIS_LOOP_737_5_VITIS_LOOP_740_6_VITIS_LOOP_fu_406.MM_OUT_2_blk_n) begin
                            if (~AESL_inst_top.MM_OUT_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_OUT_2_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_OUT_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_OUT_2_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_734_4_VITIS_LOOP_737_5_VITIS_LOOP_740_6_VITIS_LOOP_fu_406.MM_OUT_3_blk_n) begin
                            if (~AESL_inst_top.MM_OUT_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_OUT_3_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_OUT_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_OUT_3_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_734_4_VITIS_LOOP_737_5_VITIS_LOOP_740_6_VITIS_LOOP_fu_406.MM_OUT_4_blk_n) begin
                            if (~AESL_inst_top.MM_OUT_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_OUT_4_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_OUT_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_OUT_4_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_734_4_VITIS_LOOP_737_5_VITIS_LOOP_740_6_VITIS_LOOP_fu_406.MM_OUT_5_blk_n) begin
                            if (~AESL_inst_top.MM_OUT_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_OUT_5_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_OUT_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_OUT_5_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_734_4_VITIS_LOOP_737_5_VITIS_LOOP_740_6_VITIS_LOOP_fu_406.MM_OUT_6_blk_n) begin
                            if (~AESL_inst_top.MM_OUT_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_OUT_6_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_OUT_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_OUT_6_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_734_4_VITIS_LOOP_737_5_VITIS_LOOP_740_6_VITIS_LOOP_fu_406.MM_OUT_7_blk_n) begin
                            if (~AESL_inst_top.MM_OUT_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_OUT_7_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_OUT_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_OUT_7_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_734_4_VITIS_LOOP_737_5_VITIS_LOOP_740_6_VITIS_LOOP_fu_406.MM_OUT_8_blk_n) begin
                            if (~AESL_inst_top.MM_OUT_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_OUT_8_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_OUT_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_OUT_8_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_734_4_VITIS_LOOP_737_5_VITIS_LOOP_740_6_VITIS_LOOP_fu_406.MM_OUT_9_blk_n) begin
                            if (~AESL_inst_top.MM_OUT_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_OUT_9_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_OUT_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_OUT_9_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_734_4_VITIS_LOOP_737_5_VITIS_LOOP_740_6_VITIS_LOOP_fu_406.MM_OUT_10_blk_n) begin
                            if (~AESL_inst_top.MM_OUT_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_OUT_10_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_OUT_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_OUT_10_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_734_4_VITIS_LOOP_737_5_VITIS_LOOP_740_6_VITIS_LOOP_fu_406.MM_OUT_11_blk_n) begin
                            if (~AESL_inst_top.MM_OUT_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_OUT_11_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_OUT_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_OUT_11_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_734_4_VITIS_LOOP_737_5_VITIS_LOOP_740_6_VITIS_LOOP_fu_406.MM_OUT_12_blk_n) begin
                            if (~AESL_inst_top.MM_OUT_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_OUT_12_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_OUT_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_OUT_12_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_734_4_VITIS_LOOP_737_5_VITIS_LOOP_740_6_VITIS_LOOP_fu_406.MM_OUT_13_blk_n) begin
                            if (~AESL_inst_top.MM_OUT_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_OUT_13_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_OUT_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_OUT_13_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_734_4_VITIS_LOOP_737_5_VITIS_LOOP_740_6_VITIS_LOOP_fu_406.MM_OUT_14_blk_n) begin
                            if (~AESL_inst_top.MM_OUT_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_OUT_14_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_OUT_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_OUT_14_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.grp_ResOutput_Pipeline_VITIS_LOOP_734_4_VITIS_LOOP_737_5_VITIS_LOOP_740_6_VITIS_LOOP_fu_406.MM_OUT_15_blk_n) begin
                            if (~AESL_inst_top.MM_OUT_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.MM_OUT_15_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.MM_OUT_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.MM_OUT_15_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.MM_OUT_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.R_blk_n) begin
                            if (~AESL_inst_top.R_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.R_c_U' written by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.R_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.R_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.R_c_U' read by process 'top.ConvertToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.R_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    0: begin
                        if (~AESL_inst_top.ResOutput_U0.output_r_blk_n) begin
                            if (~AESL_inst_top.Output_r_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.Output_r_c_U' written by process 'top.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Output_r_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.Output_r_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.Output_r_c_U' read by process 'top.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.Output_r_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.start_for_ResOutput_U0_U.if_empty_n & AESL_inst_top.ResOutput_U0.ap_idle & ~AESL_inst_top.start_for_ResOutput_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'top.start_for_ResOutput_U0_U' written by process 'top.entry_proc_U0',");
                        end
                    end
                    5: begin
                        if (~AESL_inst_top.ResOutput_U0.C_blk_n) begin
                            if (~AESL_inst_top.C_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.C_c_U' written by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.C_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.C_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.C_c_U' read by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.C_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.P_blk_n) begin
                            if (~AESL_inst_top.P_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.P_c_U' written by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.P_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.P_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.P_c_U' read by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.P_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_top.ResOutput_U0.S_blk_n) begin
                            if (~AESL_inst_top.S_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.S_c_U' written by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.S_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.S_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.S_c_U' read by process 'top.Sliding_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.S_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    13: begin
                        if (~AESL_inst_top.ResOutput_U0.K_blk_n) begin
                            if (~AESL_inst_top.K_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'top.K_c_U' written by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.K_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_top.K_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'top.K_c_U' read by process 'top.ConvToOutStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path top.K_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
            endcase
        end
    endtask

    // report
    initial begin : report_deadlock
        integer cycle_id;
        integer cycle_comp_id;
        integer record_time;
        wait (dl_reset == 1);
        cycle_id = 1;
        record_time = 0;
        while (1) begin
            @ (negedge dl_clock);
            case (CS_fsm)
                ST_DL_DETECTED: begin
                    cycle_comp_id = 2;
                    if (dl_detect_reg != dl_done_reg) begin
                        if (dl_done_reg == 'b0) begin
                            print_dl_head;
                            record_time = $time;
                        end
                        print_cycle_start(proc_path(origin), cycle_id);
                        cycle_id = cycle_id + 1;
                    end
                    else begin
                        print_dl_end((cycle_id - 1),record_time);
                        @(negedge dl_clock);
                        @(negedge dl_clock);
                        $finish;
                    end
                end
                ST_DL_REPORT: begin
                    if ((|(dl_in_vec)) & ~(|(dl_in_vec & origin_reg))) begin
                        print_cycle_chan_comp(dl_in_vec_reg, dl_in_vec);
                        print_cycle_proc_comp(proc_path(dl_in_vec), cycle_comp_id);
                        cycle_comp_id = cycle_comp_id + 1;
                    end
                    else begin
                        print_cycle_chan_comp(dl_in_vec_reg, dl_in_vec);
                    end
                end
            endcase
        end
    end
 
endmodule
